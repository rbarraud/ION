--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Built for project 'Opcode tester'.
--------------------------------------------------------------------------------
-- This file contains object code in the form of a VHDL byte table constant.
-- This constant can be used to initialize FPGA memories for synthesis or
-- simulation.
-- Note that the object code is stored as a plain byte table in byte address
-- order. This table knows nothing of data endianess and can be used to
-- initialize 32-, 16- or 8-bit-wide memory -- memory initialization functions
-- can be found in package mips_pkg.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ION_MAIN_PKG.all;

package sim_params_pkg is

-- Hardcoded simulation parameters ---------------------------------------------

-- Simulation clock rate
constant CLOCK_RATE : integer   := 50e6;
-- Simulation clock period
constant T : time               := (1.0e9/real(CLOCK_RATE)) * 1 ns;

-- Other simulation parameters -------------------------------------------------

constant SIMULATION_LENGTH : integer := 140000;
constant LOG_TRIGGER_ADDRESS : t_word := X"bfc00000";
constant SRAM_SIZE : integer := 1024;
constant PROM_SIZE : integer := 0;
constant BRAM_SIZE : integer := 4096;


-- Memory initialization data --------------------------------------------------

constant obj_code : t_obj_code(0 to 5339) := (
  X"10", X"00", X"00", X"79", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"40", X"1a", X"68", X"00", X"00", X"1a", X"d0", X"82", 
  X"33", X"5a", X"00", X"1f", X"34", X"1b", X"00", X"08", 
  X"13", X"5b", X"00", X"09", X"23", X"7b", X"00", X"01", 
  X"13", X"5b", X"00", X"05", X"23", X"7b", X"00", X"01", 
  X"17", X"5b", X"00", X"0e", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"79", X"20", X"84", X"00", X"04", 
  X"0b", X"f0", X"00", X"79", X"20", X"84", X"00", X"05", 
  X"40", X"1a", X"68", X"00", X"00", X"1a", X"d0", X"82", 
  X"33", X"5a", X"00", X"1f", X"23", X"5a", X"ff", X"f8", 
  X"17", X"40", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"20", X"44", X"00", X"22", X"42", X"00", X"00", X"18", 
  X"34", X"04", X"00", X"99", X"0b", X"f0", X"00", X"79", 
  X"20", X"84", X"00", X"0f", X"42", X"00", X"00", X"18", 
  X"3c", X"1c", X"00", X"00", X"27", X"9c", X"7f", X"f0", 
  X"3c", X"04", X"00", X"00", X"24", X"84", X"00", X"00", 
  X"3c", X"05", X"00", X"00", X"24", X"a5", X"00", X"40", 
  X"00", X"00", X"00", X"00", X"3c", X"14", X"20", X"00", 
  X"34", X"15", X"00", X"0a", X"34", X"16", X"00", X"58", 
  X"34", X"17", X"00", X"0d", X"34", X"18", X"0f", X"80", 
  X"3c", X"1a", X"20", X"01", X"34", X"1b", X"00", X"00", 
  X"af", X"5b", X"00", X"34", X"40", X"1a", X"60", X"00", 
  X"40", X"1a", X"68", X"00", X"34", X"04", X"00", X"42", 
  X"3c", X"1a", X"00", X"40", X"37", X"5a", X"00", X"10", 
  X"40", X"9a", X"60", X"00", X"00", X"00", X"00", X"00", 
  X"34", X"04", X"00", X"34", X"40", X"1b", X"68", X"00", 
  X"00", X"00", X"00", X"00", X"40", X"1b", X"60", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"41", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"72", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"69", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"74", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"68", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"34", X"03", X"00", X"05", X"34", X"04", X"00", X"3c", 
  X"00", X"64", X"10", X"20", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"62", X"a2", X"82", X"00", X"00", 
  X"34", X"04", X"00", X"3c", X"20", X"82", X"00", X"05", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"63", 
  X"a2", X"82", X"00", X"00", X"34", X"04", X"00", X"32", 
  X"24", X"85", X"00", X"0f", X"a2", X"85", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"64", X"a2", X"82", X"00", X"00", 
  X"34", X"03", X"00", X"05", X"34", X"04", X"00", X"3c", 
  X"00", X"64", X"10", X"20", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"69", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"0a", X"34", X"03", X"00", X"0c", 
  X"00", X"43", X"20", X"2a", X"20", X"85", X"00", X"40", 
  X"a2", X"85", X"00", X"00", X"00", X"62", X"20", X"2a", 
  X"20", X"85", X"00", X"42", X"a2", X"85", X"00", X"00", 
  X"24", X"02", X"ff", X"f0", X"00", X"43", X"20", X"2a", 
  X"20", X"85", X"00", X"42", X"a2", X"85", X"00", X"00", 
  X"00", X"62", X"20", X"2a", X"20", X"85", X"00", X"44", 
  X"a2", X"85", X"00", X"00", X"24", X"03", X"ff", X"ff", 
  X"00", X"43", X"20", X"2a", X"20", X"85", X"00", X"44", 
  X"a2", X"85", X"00", X"00", X"00", X"62", X"20", X"2a", 
  X"20", X"85", X"00", X"46", X"a2", X"85", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6a", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"0a", X"28", X"44", X"00", X"0c", 
  X"20", X"85", X"00", X"40", X"a2", X"85", X"00", X"00", 
  X"28", X"44", X"00", X"08", X"20", X"85", X"00", X"42", 
  X"a2", X"85", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"6b", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"00", X"0a", 
  X"2c", X"44", X"00", X"0c", X"20", X"85", X"00", X"40", 
  X"a2", X"85", X"00", X"00", X"2c", X"44", X"00", X"08", 
  X"20", X"85", X"00", X"42", X"a2", X"85", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6c", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"0a", X"34", X"03", X"00", X"0c", 
  X"00", X"43", X"20", X"2a", X"20", X"85", X"00", X"40", 
  X"a2", X"85", X"00", X"00", X"00", X"62", X"20", X"2a", 
  X"20", X"85", X"00", X"42", X"a2", X"85", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6d", X"a2", X"82", X"00", X"00", 
  X"34", X"03", X"00", X"46", X"34", X"04", X"00", X"05", 
  X"00", X"64", X"10", X"22", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6e", X"a2", X"82", X"00", X"00", 
  X"34", X"03", X"00", X"46", X"34", X"04", X"00", X"05", 
  X"00", X"64", X"10", X"22", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"42", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"72", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"6e", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"63", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"68", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"10", X"00", X"00", X"02", X"a2", X"8a", X"00", X"00", 
  X"a2", X"96", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"62", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"0e", X"00", X"45", X"34", X"0f", X"00", X"58", 
  X"04", X"11", X"00", X"05", X"a2", X"8a", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"10", X"00", X"00", X"06", 
  X"a2", X"8e", X"00", X"00", X"a2", X"8f", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"a2", X"8c", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"63", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"02", X"00", X"64", X"34", X"03", X"00", X"7b", 
  X"34", X"04", X"00", X"7b", X"10", X"43", X"00", X"05", 
  X"a2", X"8a", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"10", X"64", X"00", X"02", X"a2", X"8c", X"00", X"00", 
  X"a2", X"96", X"00", X"00", X"a2", X"8d", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"64", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"0f", X"00", X"58", X"34", X"02", X"00", X"64", 
  X"3c", X"03", X"ff", X"ff", X"34", X"63", X"12", X"34", 
  X"34", X"04", X"00", X"7b", X"04", X"61", X"00", X"05", 
  X"a2", X"8a", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"04", X"41", X"00", X"02", X"a2", X"8c", X"00", X"00", 
  X"a2", X"96", X"00", X"00", X"04", X"01", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"a2", X"8f", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"65", 
  X"a2", X"82", X"00", X"00", X"34", X"0a", X"00", X"41", 
  X"34", X"0b", X"00", X"42", X"34", X"0c", X"00", X"43", 
  X"34", X"0d", X"00", X"44", X"34", X"0e", X"00", X"45", 
  X"34", X"0f", X"00", X"58", X"3c", X"03", X"ff", X"ff", 
  X"34", X"63", X"12", X"34", X"04", X"71", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"a2", X"8a", X"00", X"00", 
  X"04", X"11", X"00", X"05", X"00", X"00", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"10", X"00", X"00", X"06", 
  X"a2", X"8e", X"00", X"00", X"a2", X"8f", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"a2", X"8c", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"66", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"02", X"00", X"64", X"3c", X"03", X"ff", X"ff", 
  X"34", X"63", X"12", X"34", X"1c", X"60", X"00", X"05", 
  X"a2", X"8a", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"1c", X"40", X"00", X"02", X"a2", X"8c", X"00", X"00", 
  X"a2", X"96", X"00", X"00", X"a2", X"8d", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"67", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"02", X"00", X"64", X"3c", X"03", X"ff", X"ff", 
  X"34", X"63", X"12", X"34", X"18", X"40", X"00", X"05", 
  X"a2", X"8a", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"18", X"60", X"00", X"02", X"a2", X"8c", X"00", X"00", 
  X"a2", X"96", X"00", X"00", X"18", X"00", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"68", 
  X"a2", X"82", X"00", X"00", X"34", X"0a", X"00", X"41", 
  X"34", X"0b", X"00", X"42", X"34", X"0c", X"00", X"43", 
  X"34", X"0d", X"00", X"44", X"34", X"0e", X"00", X"45", 
  X"34", X"02", X"00", X"64", X"3c", X"03", X"ff", X"ff", 
  X"34", X"63", X"12", X"34", X"34", X"04", X"00", X"00", 
  X"04", X"40", X"00", X"05", X"a2", X"8a", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"04", X"60", X"00", X"02", 
  X"a2", X"8c", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"04", X"80", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"a2", X"8e", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"69", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"0e", X"00", X"45", X"34", X"0f", X"00", X"58", 
  X"3c", X"03", X"ff", X"ff", X"34", X"63", X"12", X"34", 
  X"04", X"10", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"a2", X"8a", X"00", X"00", X"04", X"70", X"00", X"05", 
  X"00", X"00", X"00", X"00", X"a2", X"8d", X"00", X"00", 
  X"10", X"00", X"00", X"06", X"a2", X"8e", X"00", X"00", 
  X"a2", X"8f", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"a2", X"8c", X"00", X"00", 
  X"a2", X"96", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"6a", 
  X"a2", X"82", X"00", X"00", X"34", X"0a", X"00", X"41", 
  X"34", X"0b", X"00", X"42", X"34", X"0c", X"00", X"43", 
  X"34", X"0d", X"00", X"44", X"34", X"02", X"00", X"64", 
  X"34", X"03", X"00", X"7b", X"34", X"04", X"00", X"7b", 
  X"14", X"64", X"00", X"05", X"a2", X"8a", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"14", X"43", X"00", X"02", 
  X"a2", X"8c", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"6b", 
  X"a2", X"82", X"00", X"00", X"34", X"0a", X"00", X"41", 
  X"34", X"0b", X"00", X"42", X"34", X"0f", X"00", X"58", 
  X"0b", X"f0", X"01", X"ed", X"a2", X"8a", X"00", X"00", 
  X"a2", X"8f", X"00", X"00", X"a2", X"8b", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6c", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"0e", X"00", X"45", X"34", X"0f", X"00", X"58", 
  X"0f", X"f0", X"01", X"fe", X"a2", X"8a", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"10", X"00", X"00", X"06", 
  X"a2", X"8e", X"00", X"00", X"a2", X"8f", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"a2", X"8c", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6d", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0c", X"00", X"43", X"34", X"0d", X"00", X"44", 
  X"34", X"0e", X"00", X"45", X"34", X"0f", X"00", X"58", 
  X"3c", X"03", X"bf", X"c0", X"24", X"63", X"08", X"50", 
  X"00", X"60", X"f8", X"09", X"a2", X"8a", X"00", X"00", 
  X"a2", X"8d", X"00", X"00", X"10", X"00", X"00", X"06", 
  X"a2", X"8e", X"00", X"00", X"a2", X"8f", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"a2", X"8c", X"00", X"00", X"a2", X"96", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"6e", X"a2", X"82", X"00", X"00", 
  X"34", X"0a", X"00", X"41", X"34", X"0b", X"00", X"42", 
  X"34", X"0f", X"00", X"58", X"3c", X"03", X"bf", X"c0", 
  X"24", X"63", X"08", X"90", X"00", X"60", X"00", X"08", 
  X"a2", X"8a", X"00", X"00", X"a2", X"8f", X"00", X"00", 
  X"a2", X"8b", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"6f", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"00", X"41", 
  X"00", X"00", X"00", X"00", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"70", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"7a", X"34", X"04", X"00", X"3b", 
  X"00", X"00", X"00", X"0d", X"20", X"84", X"00", X"01", 
  X"a2", X"84", X"00", X"00", X"00", X"00", X"00", X"0d", 
  X"80", X"42", X"00", X"10", X"00", X"00", X"00", X"0d", 
  X"0b", X"f0", X"02", X"3a", X"20", X"84", X"00", X"05", 
  X"20", X"84", X"00", X"01", X"00", X"00", X"00", X"0d", 
  X"a2", X"84", X"00", X"00", X"20", X"84", X"00", X"01", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"71", X"a2", X"82", X"00", X"00", 
  X"34", X"05", X"00", X"41", X"34", X"02", X"00", X"00", 
  X"34", X"04", X"00", X"00", X"00", X"00", X"00", X"0c", 
  X"20", X"84", X"ff", X"de", X"14", X"80", X"00", X"12", 
  X"00", X"00", X"00", X"00", X"a2", X"85", X"00", X"00", 
  X"20", X"a5", X"00", X"01", X"34", X"02", X"00", X"14", 
  X"00", X"00", X"00", X"0c", X"80", X"42", X"00", X"10", 
  X"20", X"84", X"ff", X"ca", X"14", X"80", X"00", X"0a", 
  X"00", X"00", X"00", X"00", X"a2", X"85", X"00", X"00", 
  X"20", X"05", X"00", X"01", X"00", X"00", X"00", X"0c", 
  X"0b", X"f0", X"02", X"56", X"20", X"84", X"00", X"05", 
  X"20", X"84", X"00", X"01", X"20", X"84", X"00", X"01", 
  X"0b", X"f0", X"02", X"5c", X"00", X"00", X"00", X"00", 
  X"34", X"05", X"00", X"3f", X"a2", X"85", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"4c", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"6f", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"64", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"00", X"18", X"10", X"25", X"3c", X"03", X"41", X"42", 
  X"34", X"63", X"43", X"fc", X"ac", X"43", X"00", X"10", 
  X"80", X"44", X"00", X"10", X"a2", X"84", X"00", X"00", 
  X"80", X"44", X"00", X"11", X"00", X"00", X"00", X"00", 
  X"a2", X"84", X"00", X"00", X"80", X"44", X"00", X"12", 
  X"00", X"00", X"00", X"00", X"a2", X"84", X"00", X"00", 
  X"80", X"42", X"00", X"13", X"00", X"00", X"00", X"00", 
  X"00", X"02", X"1a", X"03", X"20", X"63", X"00", X"45", 
  X"a2", X"83", X"00", X"00", X"20", X"42", X"00", X"49", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"62", 
  X"a2", X"82", X"00", X"00", X"00", X"18", X"10", X"25", 
  X"3c", X"03", X"41", X"42", X"34", X"63", X"43", X"44", 
  X"ac", X"43", X"00", X"10", X"80", X"44", X"00", X"10", 
  X"a2", X"84", X"00", X"00", X"80", X"44", X"00", X"11", 
  X"a2", X"84", X"00", X"00", X"80", X"44", X"00", X"12", 
  X"a2", X"84", X"00", X"00", X"80", X"42", X"00", X"13", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"63", 
  X"a2", X"82", X"00", X"00", X"00", X"18", X"10", X"25", 
  X"3c", X"03", X"00", X"41", X"34", X"63", X"00", X"42", 
  X"ac", X"43", X"00", X"10", X"84", X"44", X"00", X"10", 
  X"a2", X"84", X"00", X"00", X"84", X"42", X"00", X"12", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"64", 
  X"a2", X"82", X"00", X"00", X"00", X"18", X"10", X"25", 
  X"3c", X"03", X"00", X"41", X"34", X"63", X"00", X"42", 
  X"ac", X"43", X"00", X"10", X"84", X"44", X"00", X"10", 
  X"a2", X"84", X"00", X"00", X"84", X"42", X"00", X"12", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"65", 
  X"a2", X"82", X"00", X"00", X"00", X"18", X"10", X"25", 
  X"24", X"03", X"00", X"41", X"ac", X"43", X"00", X"10", 
  X"34", X"03", X"00", X"00", X"8c", X"42", X"00", X"10", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"67", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"00", X"41", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"68", 
  X"a2", X"82", X"00", X"00", X"00", X"18", X"20", X"25", 
  X"34", X"02", X"41", X"42", X"a4", X"82", X"00", X"10", 
  X"80", X"83", X"00", X"10", X"a2", X"83", X"00", X"00", 
  X"80", X"82", X"00", X"11", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"69", X"a2", X"82", X"00", X"00", 
  X"00", X"18", X"10", X"25", X"3c", X"03", X"41", X"42", 
  X"34", X"63", X"43", X"44", X"ac", X"43", X"00", X"10", 
  X"80", X"44", X"00", X"10", X"a2", X"84", X"00", X"00", 
  X"80", X"44", X"00", X"11", X"a2", X"84", X"00", X"00", 
  X"80", X"44", X"00", X"12", X"a2", X"84", X"00", X"00", 
  X"80", X"42", X"00", X"13", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"4c", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"6f", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"67", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"69", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"63", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"07", X"41", X"34", X"03", X"60", X"f3", 
  X"00", X"43", X"20", X"24", X"a2", X"84", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"62", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"07", X"41", X"30", X"44", X"60", X"f3", 
  X"a2", X"84", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"63", 
  X"a2", X"82", X"00", X"00", X"3c", X"02", X"00", X"41", 
  X"00", X"02", X"1c", X"02", X"a2", X"83", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"64", X"a2", X"82", X"00", X"00", 
  X"3c", X"02", X"f0", X"ff", X"34", X"42", X"f0", X"8e", 
  X"3c", X"03", X"0f", X"0f", X"34", X"63", X"0f", X"30", 
  X"00", X"43", X"20", X"27", X"a2", X"84", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"65", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"40", X"34", X"03", X"00", X"01", 
  X"00", X"43", X"20", X"25", X"a2", X"84", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"66", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"40", X"34", X"44", X"00", X"01", 
  X"a2", X"84", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"67", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"f0", X"43", 
  X"34", X"03", X"f0", X"02", X"00", X"43", X"20", X"26", 
  X"a2", X"84", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"68", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"f0", X"43", 
  X"38", X"44", X"f0", X"02", X"a2", X"84", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"4d", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"6f", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"76", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"65", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"53", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"68", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"69", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"66", X"a2", X"82", X"00", X"00", 
  X"34", X"02", X"00", X"74", X"a2", X"82", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"61", X"a2", X"82", X"00", X"00", 
  X"3c", X"02", X"40", X"41", X"34", X"42", X"42", X"43", 
  X"00", X"02", X"1a", X"00", X"00", X"03", X"1e", X"02", 
  X"a2", X"83", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"62", 
  X"a2", X"82", X"00", X"00", X"3c", X"02", X"40", X"41", 
  X"34", X"42", X"42", X"43", X"34", X"03", X"00", X"08", 
  X"00", X"62", X"18", X"04", X"00", X"03", X"1e", X"02", 
  X"a2", X"83", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"63", 
  X"a2", X"82", X"00", X"00", X"3c", X"02", X"40", X"41", 
  X"34", X"42", X"42", X"43", X"00", X"02", X"1c", X"03", 
  X"a2", X"83", X"00", X"00", X"3c", X"02", X"84", X"00", 
  X"00", X"02", X"1e", X"43", X"20", X"63", X"ff", X"80", 
  X"a2", X"83", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"64", 
  X"a2", X"82", X"00", X"00", X"3c", X"02", X"40", X"41", 
  X"34", X"42", X"42", X"43", X"34", X"03", X"00", X"10", 
  X"00", X"62", X"18", X"07", X"a2", X"83", X"00", X"00", 
  X"34", X"03", X"00", X"19", X"3c", X"02", X"84", X"00", 
  X"00", X"62", X"18", X"07", X"20", X"63", X"ff", X"80", 
  X"a2", X"83", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"65", 
  X"a2", X"82", X"00", X"00", X"3c", X"02", X"40", X"41", 
  X"34", X"42", X"42", X"43", X"00", X"02", X"1c", X"02", 
  X"a2", X"83", X"00", X"00", X"3c", X"02", X"84", X"00", 
  X"00", X"02", X"1e", X"42", X"a2", X"83", X"00", X"00", 
  X"a2", X"97", X"00", X"00", X"a2", X"95", X"00", X"00", 
  X"34", X"02", X"00", X"66", X"a2", X"82", X"00", X"00", 
  X"3c", X"02", X"40", X"41", X"34", X"42", X"42", X"43", 
  X"34", X"03", X"00", X"10", X"00", X"62", X"20", X"06", 
  X"a2", X"84", X"00", X"00", X"34", X"03", X"00", X"19", 
  X"3c", X"02", X"84", X"00", X"00", X"62", X"18", X"06", 
  X"a2", X"83", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"02", X"00", X"44", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"00", X"6f", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"00", X"6e", 
  X"a2", X"82", X"00", X"00", X"34", X"02", X"00", X"65", 
  X"a2", X"82", X"00", X"00", X"a2", X"97", X"00", X"00", 
  X"a2", X"95", X"00", X"00", X"34", X"10", X"a5", X"a5", 
  X"34", X"11", X"00", X"0f", X"34", X"12", X"00", X"01", 
  X"24", X"13", X"ff", X"ff", X"24", X"14", X"fc", X"18", 
  X"3c", X"15", X"80", X"00", X"3c", X"16", X"7f", X"ff", 
  X"36", X"d6", X"ff", X"ff", X"02", X"00", X"40", X"21", 
  X"02", X"20", X"48", X"21", X"01", X"31", X"40", X"20", 
  X"02", X"00", X"40", X"21", X"02", X"20", X"48", X"21", 
  X"01", X"33", X"40", X"20", X"02", X"00", X"40", X"21", 
  X"02", X"20", X"48", X"21", X"01", X"34", X"40", X"20", 
  X"02", X"00", X"40", X"21", X"02", X"c0", X"48", X"21", 
  X"01", X"36", X"40", X"20", X"02", X"00", X"40", X"21", 
  X"02", X"a0", X"48", X"21", X"01", X"35", X"40", X"20", 
  X"02", X"00", X"40", X"21", X"02", X"a0", X"48", X"21", 
  X"21", X"28", X"ff", X"ff", X"02", X"00", X"40", X"21", 
  X"02", X"a0", X"48", X"21", X"21", X"28", X"00", X"0f", 
  X"02", X"00", X"40", X"21", X"02", X"60", X"48", X"21", 
  X"21", X"28", X"00", X"02", X"02", X"00", X"40", X"21", 
  X"02", X"20", X"48", X"21", X"21", X"28", X"00", X"02", 
  X"02", X"00", X"40", X"21", X"02", X"c0", X"48", X"21", 
  X"21", X"28", X"00", X"02", X"02", X"00", X"40", X"21", 
  X"02", X"a0", X"48", X"21", X"25", X"28", X"ff", X"ff", 
  X"02", X"00", X"40", X"21", X"02", X"a0", X"48", X"21", 
  X"25", X"28", X"00", X"0f", X"02", X"00", X"40", X"21", 
  X"02", X"60", X"48", X"21", X"25", X"28", X"00", X"02", 
  X"02", X"00", X"40", X"21", X"02", X"20", X"48", X"21", 
  X"25", X"28", X"00", X"02", X"02", X"00", X"40", X"21", 
  X"02", X"c0", X"48", X"21", X"25", X"28", X"00", X"02", 
  X"02", X"00", X"40", X"21", X"02", X"20", X"48", X"21", 
  X"01", X"31", X"40", X"21", X"02", X"00", X"40", X"21", 
  X"02", X"20", X"48", X"21", X"01", X"33", X"40", X"21", 
  X"02", X"00", X"40", X"21", X"02", X"20", X"48", X"21", 
  X"01", X"34", X"40", X"21", X"02", X"00", X"40", X"21", 
  X"02", X"c0", X"48", X"21", X"01", X"36", X"40", X"21", 
  X"02", X"00", X"40", X"21", X"02", X"a0", X"48", X"21", 
  X"01", X"35", X"40", X"21", X"02", X"00", X"40", X"21", 
  X"02", X"40", X"48", X"21", X"01", X"31", X"40", X"22", 
  X"02", X"00", X"40", X"21", X"02", X"20", X"48", X"21", 
  X"01", X"33", X"40", X"20", X"02", X"00", X"40", X"21", 
  X"02", X"20", X"48", X"21", X"01", X"34", X"40", X"20", 
  X"02", X"00", X"40", X"21", X"02", X"c0", X"48", X"21", 
  X"01", X"36", X"40", X"20", X"02", X"00", X"40", X"21", 
  X"02", X"a0", X"48", X"21", X"01", X"35", X"40", X"20", 
  X"34", X"06", X"a5", X"a5", X"34", X"04", X"00", X"0f", 
  X"34", X"05", X"00", X"01", X"00", X"e0", X"10", X"21", 
  X"00", X"85", X"10", X"2a", X"00", X"e0", X"10", X"21", 
  X"00", X"a4", X"10", X"2a", X"00", X"e0", X"10", X"21", 
  X"28", X"82", X"00", X"01", X"00", X"e0", X"10", X"21", 
  X"28", X"a2", X"00", X"0f", X"00", X"e0", X"10", X"21", 
  X"2c", X"82", X"00", X"01", X"00", X"e0", X"10", X"21", 
  X"2c", X"a2", X"00", X"0f", X"34", X"05", X"a5", X"a5", 
  X"24", X"04", X"04", X"05", X"24", X"84", X"f8", X"30", 
  X"2c", X"85", X"03", X"e8", X"3c", X"10", X"7f", X"ff", 
  X"36", X"10", X"ff", X"ff", X"36", X"31", X"03", X"e8", 
  X"36", X"31", X"00", X"0f", X"36", X"31", X"00", X"02", 
  X"3c", X"14", X"80", X"00", X"24", X"15", X"fc", X"17", 
  X"24", X"16", X"ff", X"f0", X"24", X"17", X"ff", X"fd", 
  X"1e", X"20", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"34", X"42", X"55", X"00", X"1e", X"e0", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"34", X"42", X"55", X"01", 
  X"1e", X"00", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"34", X"42", X"55", X"02", X"1e", X"80", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"34", X"42", X"55", X"03", 
  X"06", X"21", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"34", X"42", X"55", X"00", X"06", X"e1", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"34", X"42", X"55", X"01", 
  X"06", X"01", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"34", X"42", X"55", X"02", X"06", X"81", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"34", X"42", X"55", X"03", 
  X"06", X"20", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"34", X"42", X"55", X"00", X"06", X"e0", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"34", X"42", X"55", X"01", 
  X"06", X"00", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"34", X"42", X"55", X"02", X"06", X"80", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"34", X"42", X"55", X"03", 
  X"0b", X"f0", X"04", X"14", X"00", X"00", X"00", X"00", 
  X"3c", X"04", X"00", X"01", X"40", X"84", X"60", X"00", 
  X"3c", X"04", X"00", X"00", X"24", X"84", X"00", X"00", 
  X"24", X"06", X"00", X"00", X"24", X"05", X"00", X"ff", 
  X"ac", X"86", X"00", X"00", X"00", X"c5", X"08", X"2a", 
  X"14", X"20", X"ff", X"fd", X"20", X"c6", X"00", X"01", 
  X"24", X"04", X"00", X"00", X"24", X"06", X"00", X"00", 
  X"24", X"05", X"00", X"ff", X"8c", X"80", X"00", X"00", 
  X"20", X"84", X"00", X"10", X"00", X"c5", X"08", X"2a", 
  X"14", X"20", X"ff", X"fc", X"20", X"c6", X"00", X"01", 
  X"3c", X"05", X"00", X"02", X"34", X"a5", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"40", X"85", X"60", X"00", 
  X"3c", X"1b", X"00", X"00", X"27", X"7b", X"00", X"3c", 
  X"af", X"7d", X"ff", X"f0", X"af", X"7f", X"ff", X"ec", 
  X"af", X"68", X"ff", X"e8", X"af", X"69", X"ff", X"e4", 
  X"af", X"6a", X"ff", X"e0", X"03", X"60", X"e8", X"21", 
  X"40", X"08", X"70", X"00", X"8d", X"1a", X"00", X"00", 
  X"40", X"1b", X"68", X"00", X"07", X"70", X"00", X"2d", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"4e", X"82", 
  X"39", X"28", X"00", X"1f", X"11", X"00", X"00", X"1f", 
  X"39", X"28", X"00", X"1c", X"11", X"00", X"00", X"13", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"8f", X"aa", X"ff", X"e0", 
  X"8f", X"a9", X"ff", X"e4", X"8f", X"a8", X"ff", X"e8", 
  X"8f", X"bf", X"ff", X"ec", X"8f", X"bd", X"ff", X"f0", 
  X"40", X"1b", X"70", X"00", X"40", X"1a", X"68", X"00", 
  X"00", X"1a", X"d7", X"c2", X"33", X"5a", X"00", X"01", 
  X"17", X"40", X"00", X"03", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"42", X"00", X"00", X"10", X"33", X"5b", X"00", X"3f", 
  X"3b", X"68", X"00", X"20", X"11", X"00", X"00", X"14", 
  X"3b", X"68", X"00", X"21", X"11", X"00", X"00", X"1c", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"0b", X"f0", X"04", X"41", 
  X"00", X"00", X"00", X"00", X"33", X"5b", X"00", X"3f", 
  X"3b", X"68", X"00", X"00", X"11", X"00", X"00", X"1e", 
  X"3b", X"68", X"00", X"04", X"11", X"00", X"00", X"29", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"0b", X"f0", X"04", X"41", 
  X"00", X"00", X"00", X"00", X"8d", X"1a", X"00", X"04", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"0f", X"f0", X"04", X"eb", X"3c", X"0a", X"80", X"00", 
  X"00", X"00", X"40", X"21", X"03", X"6a", X"48", X"24", 
  X"15", X"20", X"00", X"03", X"00", X"0a", X"50", X"42", 
  X"15", X"40", X"ff", X"fc", X"25", X"08", X"00", X"01", 
  X"0b", X"f0", X"04", X"a1", X"01", X"00", X"d8", X"21", 
  X"0f", X"f0", X"04", X"eb", X"3c", X"0a", X"80", X"00", 
  X"00", X"00", X"40", X"21", X"03", X"6a", X"48", X"24", 
  X"11", X"20", X"00", X"03", X"00", X"0a", X"50", X"42", 
  X"15", X"40", X"ff", X"fc", X"25", X"08", X"00", X"01", 
  X"0b", X"f0", X"04", X"a1", X"01", X"00", X"d8", X"21", 
  X"0f", X"f0", X"04", X"eb", X"00", X"00", X"00", X"00", 
  X"00", X"1a", X"41", X"82", X"31", X"08", X"00", X"1f", 
  X"00", X"1a", X"4a", X"c2", X"31", X"29", X"00", X"1f", 
  X"01", X"09", X"50", X"21", X"00", X"0a", X"50", X"23", 
  X"25", X"4a", X"00", X"1f", X"01", X"5b", X"d8", X"04", 
  X"01", X"5b", X"d8", X"06", X"0b", X"f0", X"04", X"a1", 
  X"01", X"1b", X"d8", X"06", X"0f", X"f0", X"04", X"eb", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"41", X"82", 
  X"31", X"08", X"00", X"1f", X"00", X"1a", X"4a", X"c2", 
  X"31", X"29", X"00", X"1f", X"01", X"28", X"48", X"23", 
  X"00", X"09", X"58", X"23", X"25", X"6b", X"00", X"1f", 
  X"01", X"1b", X"48", X"04", X"3c", X"0a", X"ff", X"ff", 
  X"35", X"4a", X"ff", X"ff", X"01", X"6a", X"50", X"04", 
  X"01", X"6a", X"50", X"06", X"01", X"0a", X"50", X"04", 
  X"01", X"2a", X"48", X"24", X"01", X"40", X"50", X"27", 
  X"0f", X"f0", X"04", X"eb", X"00", X"1a", X"d1", X"40", 
  X"00", X"1a", X"d1", X"42", X"03", X"6a", X"d8", X"24", 
  X"03", X"69", X"d8", X"25", X"0b", X"f0", X"04", X"a1", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"4c", X"02", 
  X"31", X"29", X"00", X"1f", X"3c", X"08", X"bf", X"c0", 
  X"25", X"08", X"12", X"ac", X"00", X"09", X"48", X"c0", 
  X"01", X"09", X"40", X"20", X"01", X"00", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"04", X"41", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"60", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"61", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"62", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"63", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"64", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"65", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"66", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"67", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"af", X"bb", X"ff", X"e8", X"0b", X"f0", X"04", X"a9", 
  X"af", X"bb", X"ff", X"e4", X"0b", X"f0", X"04", X"a9", 
  X"af", X"bb", X"ff", X"e0", X"0b", X"f0", X"04", X"a9", 
  X"37", X"6b", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"6c", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"6d", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"6e", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"6f", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"70", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"71", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"72", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"73", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"74", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"75", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"76", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"77", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"78", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"79", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"7a", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"7b", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"37", X"7c", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"af", X"bb", X"ff", X"ec", X"0b", X"f0", X"04", X"a9", 
  X"37", X"7e", X"00", X"00", X"0b", X"f0", X"04", X"a9", 
  X"af", X"bb", X"ff", X"f0", X"af", X"bf", X"00", X"00", 
  X"00", X"1a", X"dd", X"42", X"33", X"7b", X"00", X"1f", 
  X"3c", X"08", X"bf", X"c0", X"25", X"08", X"13", X"dc", 
  X"00", X"1b", X"d8", X"c0", X"01", X"1b", X"40", X"20", 
  X"01", X"00", X"f8", X"09", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e8", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e4", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e0", X"03", X"e0", X"00", X"08", 
  X"35", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"9a", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"f0", X"03", X"e0", X"00", X"08", 
  X"37", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"ec" );

constant sram_init : t_obj_code(0 to 0) := (others => X"00");
constant prom_init : t_obj_code(0 to 0) := (others => X"00");


end package sim_params_pkg;
