--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Built for project 'LibC Test'.
--------------------------------------------------------------------------------
-- This file contains object code in the form of a VHDL byte table constant.
-- This constant can be used to initialize FPGA memories for synthesis or
-- simulation.
-- Note that the object code is stored as a plain byte table in byte address
-- order. This table knows nothing of data endianess and can be used to
-- initialize 32-, 16- or 8-bit-wide memory -- memory initialization functions
-- can be found in package mips_pkg.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ION_MAIN_PKG.all;

package OBJ_CODE_PKG is

-- Simulation or synthesis parameters ------------------------------------------

constant CODE_MEM_SIZE : integer := 32768;
constant DATA_MEM_SIZE : integer := 32768;


-- Memory initialization data --------------------------------------------------

constant OBJ_CODE : t_obj_code(0 to 26039) := (
  X"10", X"00", X"00", X"7c", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"40", X"1a", X"68", X"00", X"00", X"1a", X"d0", X"82", 
  X"33", X"5a", X"00", X"1f", X"34", X"1b", X"00", X"08", 
  X"13", X"5b", X"00", X"09", X"23", X"7b", X"00", X"01", 
  X"13", X"5b", X"00", X"05", X"23", X"7b", X"00", X"01", 
  X"17", X"5b", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"be", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"40", X"1b", X"70", X"00", X"40", X"1a", X"68", X"00", 
  X"00", X"1a", X"d7", X"c2", X"33", X"5a", X"00", X"01", 
  X"17", X"40", X"00", X"03", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"42", X"00", X"00", X"10", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"fe", X"40", X"84", X"60", X"00", 
  X"3c", X"04", X"bf", X"c0", X"24", X"84", X"02", X"78", 
  X"00", X"80", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"3c", X"05", X"00", X"01", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"ff", X"00", X"85", X"28", X"25", 
  X"40", X"85", X"60", X"00", X"24", X"04", X"00", X"00", 
  X"24", X"06", X"00", X"00", X"24", X"05", X"00", X"ff", 
  X"ac", X"86", X"00", X"00", X"00", X"c5", X"08", X"2a", 
  X"14", X"20", X"ff", X"fd", X"20", X"c6", X"00", X"01", 
  X"24", X"04", X"00", X"00", X"24", X"06", X"00", X"00", 
  X"24", X"05", X"00", X"ff", X"8c", X"80", X"00", X"00", 
  X"20", X"84", X"00", X"10", X"00", X"c5", X"08", X"2a", 
  X"14", X"20", X"ff", X"fc", X"20", X"c6", X"00", X"01", 
  X"3c", X"05", X"00", X"02", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"ff", X"00", X"85", X"28", X"25", 
  X"03", X"e0", X"00", X"08", X"40", X"85", X"60", X"00", 
  X"3c", X"1c", X"00", X"00", X"27", X"9c", X"7f", X"f0", 
  X"3c", X"05", X"00", X"00", X"24", X"a5", X"08", X"b0", 
  X"3c", X"04", X"00", X"00", X"24", X"84", X"08", X"f4", 
  X"3c", X"1d", X"00", X"00", X"27", X"bd", X"0c", X"e8", 
  X"ac", X"a0", X"00", X"00", X"00", X"a4", X"18", X"2a", 
  X"14", X"60", X"ff", X"fd", X"24", X"a5", X"00", X"04", 
  X"3c", X"04", X"00", X"00", X"24", X"84", X"00", X"00", 
  X"3c", X"05", X"bf", X"c0", X"24", X"a5", X"5d", X"08", 
  X"10", X"a4", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"3c", X"10", X"00", X"00", X"26", X"10", X"08", X"98", 
  X"12", X"00", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"8c", X"a8", X"00", X"00", X"24", X"a5", X"00", X"04", 
  X"ac", X"88", X"00", X"00", X"24", X"84", X"00", X"04", 
  X"1e", X"00", X"ff", X"fb", X"26", X"10", X"ff", X"fc", 
  X"0f", X"f0", X"16", X"fd", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"bc", X"00", X"00", X"00", X"00", 
  X"3c", X"1b", X"00", X"00", X"27", X"7b", X"0d", X"3c", 
  X"af", X"7d", X"ff", X"f0", X"af", X"7f", X"ff", X"ec", 
  X"af", X"68", X"ff", X"e8", X"af", X"69", X"ff", X"e4", 
  X"af", X"6a", X"ff", X"e0", X"03", X"60", X"e8", X"21", 
  X"40", X"08", X"70", X"00", X"8d", X"1a", X"00", X"00", 
  X"40", X"1b", X"68", X"00", X"07", X"70", X"00", X"2d", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"4e", X"82", 
  X"39", X"28", X"00", X"1f", X"11", X"00", X"00", X"1f", 
  X"39", X"28", X"00", X"1c", X"11", X"00", X"00", X"13", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"8f", X"aa", X"ff", X"e0", 
  X"8f", X"a9", X"ff", X"e4", X"8f", X"a8", X"ff", X"e8", 
  X"8f", X"bf", X"ff", X"ec", X"8f", X"bd", X"ff", X"f0", 
  X"40", X"1b", X"70", X"00", X"40", X"1a", X"68", X"00", 
  X"00", X"1a", X"d7", X"c2", X"33", X"5a", X"00", X"01", 
  X"17", X"40", X"00", X"03", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"42", X"00", X"00", X"10", X"33", X"5b", X"00", X"3f", 
  X"3b", X"68", X"00", X"20", X"11", X"00", X"00", X"14", 
  X"3b", X"68", X"00", X"21", X"11", X"00", X"00", X"1c", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"0b", X"f0", X"00", X"d3", 
  X"00", X"00", X"00", X"00", X"33", X"5b", X"00", X"3f", 
  X"3b", X"68", X"00", X"00", X"11", X"00", X"00", X"1e", 
  X"3b", X"68", X"00", X"04", X"11", X"00", X"00", X"29", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"0b", X"f0", X"00", X"d3", 
  X"00", X"00", X"00", X"00", X"8d", X"1a", X"00", X"04", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"0f", X"f0", X"01", X"7d", X"3c", X"0a", X"80", X"00", 
  X"00", X"00", X"40", X"21", X"03", X"6a", X"48", X"24", 
  X"15", X"20", X"00", X"03", X"00", X"0a", X"50", X"42", 
  X"15", X"40", X"ff", X"fc", X"25", X"08", X"00", X"01", 
  X"0b", X"f0", X"01", X"33", X"01", X"00", X"d8", X"21", 
  X"0f", X"f0", X"01", X"7d", X"3c", X"0a", X"80", X"00", 
  X"00", X"00", X"40", X"21", X"03", X"6a", X"48", X"24", 
  X"11", X"20", X"00", X"03", X"00", X"0a", X"50", X"42", 
  X"15", X"40", X"ff", X"fc", X"25", X"08", X"00", X"01", 
  X"0b", X"f0", X"01", X"33", X"01", X"00", X"d8", X"21", 
  X"0f", X"f0", X"01", X"7d", X"00", X"00", X"00", X"00", 
  X"00", X"1a", X"41", X"82", X"31", X"08", X"00", X"1f", 
  X"00", X"1a", X"4a", X"c2", X"31", X"29", X"00", X"1f", 
  X"01", X"09", X"50", X"21", X"00", X"0a", X"50", X"23", 
  X"25", X"4a", X"00", X"1f", X"01", X"5b", X"d8", X"04", 
  X"01", X"5b", X"d8", X"06", X"0b", X"f0", X"01", X"33", 
  X"01", X"1b", X"d8", X"06", X"0f", X"f0", X"01", X"7d", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"41", X"82", 
  X"31", X"08", X"00", X"1f", X"00", X"1a", X"4a", X"c2", 
  X"31", X"29", X"00", X"1f", X"01", X"28", X"48", X"23", 
  X"00", X"09", X"58", X"23", X"25", X"6b", X"00", X"1f", 
  X"01", X"1b", X"48", X"04", X"3c", X"0a", X"ff", X"ff", 
  X"35", X"4a", X"ff", X"ff", X"01", X"6a", X"50", X"04", 
  X"01", X"6a", X"50", X"06", X"01", X"0a", X"50", X"04", 
  X"01", X"2a", X"48", X"24", X"01", X"40", X"50", X"27", 
  X"0f", X"f0", X"01", X"7d", X"00", X"1a", X"d1", X"40", 
  X"00", X"1a", X"d1", X"42", X"03", X"6a", X"d8", X"24", 
  X"03", X"69", X"d8", X"25", X"0b", X"f0", X"01", X"33", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"4c", X"02", 
  X"31", X"29", X"00", X"1f", X"3c", X"08", X"bf", X"c0", 
  X"25", X"08", X"04", X"f4", X"00", X"09", X"48", X"c0", 
  X"01", X"09", X"40", X"20", X"01", X"00", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"00", X"d3", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"60", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"61", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"62", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"63", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"64", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"65", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"66", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"67", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"af", X"bb", X"ff", X"e8", X"0b", X"f0", X"01", X"3b", 
  X"af", X"bb", X"ff", X"e4", X"0b", X"f0", X"01", X"3b", 
  X"af", X"bb", X"ff", X"e0", X"0b", X"f0", X"01", X"3b", 
  X"37", X"6b", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"6c", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"6d", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"6e", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"6f", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"70", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"71", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"72", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"73", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"74", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"75", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"76", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"77", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"78", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"79", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"7a", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"7b", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"37", X"7c", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"af", X"bb", X"ff", X"ec", X"0b", X"f0", X"01", X"3b", 
  X"37", X"7e", X"00", X"00", X"0b", X"f0", X"01", X"3b", 
  X"af", X"bb", X"ff", X"f0", X"af", X"bf", X"00", X"00", 
  X"00", X"1a", X"dd", X"42", X"33", X"7b", X"00", X"1f", 
  X"3c", X"08", X"bf", X"c0", X"25", X"08", X"06", X"24", 
  X"00", X"1b", X"d8", X"c0", X"01", X"1b", X"40", X"20", 
  X"01", X"00", X"f8", X"09", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e8", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e4", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e0", X"03", X"e0", X"00", X"08", 
  X"35", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"9a", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"f0", X"03", X"e0", X"00", X"08", 
  X"37", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"ec", X"8c", X"85", X"00", X"00", 
  X"8c", X"86", X"00", X"10", X"8c", X"83", X"00", X"14", 
  X"2c", X"a7", X"00", X"02", X"14", X"e0", X"00", X"3f", 
  X"8c", X"88", X"00", X"04", X"24", X"02", X"00", X"04", 
  X"10", X"a2", X"00", X"25", X"00", X"08", X"17", X"c0", 
  X"24", X"02", X"00", X"02", X"10", X"a2", X"00", X"3f", 
  X"00", X"08", X"17", X"c0", X"00", X"c3", X"10", X"25", 
  X"10", X"40", X"00", X"1c", X"00", X"00", X"10", X"21", 
  X"8c", X"82", X"00", X"08", X"28", X"44", X"fc", X"02", 
  X"14", X"80", X"00", X"1f", X"24", X"04", X"fc", X"02", 
  X"28", X"44", X"04", X"00", X"10", X"80", X"00", X"17", 
  X"30", X"65", X"00", X"ff", X"24", X"04", X"00", X"80", 
  X"10", X"a4", X"00", X"3c", X"24", X"64", X"00", X"7f", 
  X"00", X"83", X"18", X"2b", X"00", X"66", X"30", X"21", 
  X"00", X"80", X"18", X"21", X"3c", X"04", X"20", X"00", 
  X"00", X"c4", X"20", X"2b", X"10", X"80", X"00", X"30", 
  X"00", X"06", X"2f", X"c0", X"24", X"42", X"03", X"ff", 
  X"7c", X"c4", X"9a", X"00", X"00", X"08", X"47", X"c0", 
  X"00", X"06", X"36", X"00", X"00", X"88", X"40", X"25", 
  X"00", X"03", X"1a", X"02", X"00", X"02", X"15", X"00", 
  X"01", X"02", X"10", X"25", X"03", X"e0", X"00", X"08", 
  X"00", X"c3", X"18", X"25", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"18", X"21", X"00", X"08", X"17", X"c0", 
  X"3c", X"03", X"7f", X"f0", X"00", X"43", X"10", X"25", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"18", X"21", 
  X"00", X"82", X"10", X"23", X"28", X"44", X"00", X"39", 
  X"10", X"80", X"00", X"18", X"00", X"02", X"20", X"27", 
  X"00", X"06", X"28", X"40", X"00", X"85", X"28", X"04", 
  X"00", X"43", X"18", X"06", X"30", X"44", X"00", X"20", 
  X"00", X"a3", X"18", X"25", X"00", X"46", X"10", X"06", 
  X"00", X"44", X"18", X"0b", X"00", X"04", X"10", X"0b", 
  X"00", X"02", X"26", X"00", X"00", X"03", X"1a", X"02", 
  X"7c", X"42", X"9a", X"00", X"00", X"83", X"18", X"25", 
  X"00", X"08", X"47", X"c0", X"03", X"e0", X"00", X"08", 
  X"00", X"48", X"10", X"25", X"7c", X"c6", X"98", X"00", 
  X"3c", X"02", X"7f", X"f8", X"00", X"c2", X"10", X"25", 
  X"00", X"08", X"47", X"c0", X"03", X"e0", X"00", X"08", 
  X"00", X"48", X"10", X"25", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"18", X"21", X"00", X"00", X"10", X"21", 
  X"0b", X"f0", X"02", X"0a", X"00", X"00", X"18", X"21", 
  X"00", X"03", X"20", X"42", X"00", X"a4", X"18", X"25", 
  X"00", X"06", X"30", X"42", X"0b", X"f0", X"01", X"ea", 
  X"24", X"42", X"04", X"00", X"30", X"64", X"01", X"00", 
  X"10", X"80", X"ff", X"c7", X"3c", X"04", X"20", X"00", 
  X"24", X"64", X"00", X"80", X"00", X"83", X"18", X"2b", 
  X"00", X"66", X"30", X"21", X"0b", X"f0", X"01", X"e5", 
  X"00", X"80", X"18", X"21", X"8c", X"86", X"00", X"00", 
  X"8c", X"83", X"00", X"04", X"00", X"06", X"3f", X"c2", 
  X"7c", X"c4", X"55", X"00", X"7c", X"c2", X"98", X"00", 
  X"14", X"80", X"00", X"17", X"ac", X"a7", X"00", X"04", 
  X"00", X"43", X"20", X"25", X"10", X"80", X"00", X"23", 
  X"00", X"03", X"26", X"02", X"00", X"02", X"12", X"00", 
  X"00", X"82", X"10", X"25", X"24", X"04", X"00", X"03", 
  X"ac", X"a4", X"00", X"00", X"00", X"03", X"1a", X"00", 
  X"24", X"04", X"fc", X"01", X"3c", X"08", X"10", X"00", 
  X"00", X"03", X"37", X"c2", X"00", X"02", X"10", X"40", 
  X"00", X"c2", X"10", X"25", X"00", X"48", X"30", X"2b", 
  X"00", X"80", X"38", X"21", X"00", X"03", X"18", X"40", 
  X"14", X"c0", X"ff", X"f9", X"24", X"84", X"ff", X"ff", 
  X"ac", X"a7", X"00", X"08", X"ac", X"a2", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"ac", X"a3", X"00", X"14", 
  X"24", X"07", X"07", X"ff", X"10", X"87", X"00", X"10", 
  X"24", X"84", X"fc", X"01", X"00", X"03", X"36", X"02", 
  X"00", X"02", X"12", X"00", X"00", X"c2", X"10", X"25", 
  X"ac", X"a4", X"00", X"08", X"3c", X"06", X"10", X"00", 
  X"24", X"04", X"00", X"03", X"00", X"03", X"1a", X"00", 
  X"00", X"46", X"10", X"25", X"ac", X"a4", X"00", X"00", 
  X"ac", X"a2", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"ac", X"a3", X"00", X"14", X"24", X"02", X"00", X"02", 
  X"03", X"e0", X"00", X"08", X"ac", X"a2", X"00", X"00", 
  X"00", X"43", X"20", X"25", X"10", X"80", X"00", X"05", 
  X"7c", X"c6", X"04", X"c0", X"14", X"c0", X"00", X"06", 
  X"24", X"04", X"00", X"01", X"0b", X"f0", X"02", X"4e", 
  X"ac", X"a0", X"00", X"00", X"24", X"02", X"00", X"04", 
  X"03", X"e0", X"00", X"08", X"ac", X"a2", X"00", X"00", 
  X"0b", X"f0", X"02", X"4e", X"ac", X"a4", X"00", X"00", 
  X"8c", X"82", X"00", X"00", X"2c", X"43", X"00", X"02", 
  X"14", X"60", X"00", X"13", X"00", X"00", X"00", X"00", 
  X"8c", X"a3", X"00", X"00", X"2c", X"66", X"00", X"02", 
  X"14", X"c0", X"00", X"0f", X"24", X"06", X"00", X"04", 
  X"10", X"46", X"00", X"0f", X"00", X"00", X"00", X"00", 
  X"10", X"66", X"00", X"16", X"24", X"06", X"00", X"02", 
  X"10", X"46", X"00", X"12", X"00", X"00", X"00", X"00", 
  X"10", X"66", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"8c", X"82", X"00", X"04", X"8c", X"a3", X"00", X"04", 
  X"10", X"43", X"00", X"13", X"00", X"00", X"00", X"00", 
  X"14", X"40", X"00", X"0f", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"00", X"01", 
  X"10", X"62", X"00", X"26", X"00", X"00", X"00", X"00", 
  X"8c", X"83", X"00", X"04", X"14", X"60", X"00", X"08", 
  X"24", X"02", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"10", X"62", X"00", X"27", 
  X"00", X"00", X"00", X"00", X"8c", X"a2", X"00", X"04", 
  X"14", X"40", X"ff", X"f3", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"ff", X"ff", 
  X"8c", X"86", X"00", X"08", X"8c", X"a3", X"00", X"08", 
  X"00", X"66", X"38", X"2a", X"14", X"e0", X"ff", X"ea", 
  X"00", X"c3", X"18", X"2a", X"14", X"60", X"00", X"0f", 
  X"00", X"00", X"00", X"00", X"8c", X"a6", X"00", X"10", 
  X"8c", X"83", X"00", X"10", X"8c", X"87", X"00", X"14", 
  X"00", X"c3", X"20", X"2b", X"14", X"80", X"ff", X"e2", 
  X"8c", X"a5", X"00", X"14", X"14", X"66", X"00", X"05", 
  X"00", X"66", X"20", X"2b", X"00", X"a7", X"20", X"2b", 
  X"14", X"80", X"ff", X"dd", X"00", X"00", X"00", X"00", 
  X"00", X"66", X"20", X"2b", X"10", X"80", X"00", X"09", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"ff", X"e8", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"02", X"76", 
  X"00", X"00", X"00", X"00", X"8c", X"a3", X"00", X"04", 
  X"8c", X"82", X"00", X"04", X"03", X"e0", X"00", X"08", 
  X"00", X"62", X"10", X"23", X"14", X"c3", X"00", X"03", 
  X"00", X"e5", X"28", X"2b", X"14", X"a0", X"ff", X"f5", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"10", X"21", X"8c", X"83", X"00", X"00", 
  X"2c", X"62", X"00", X"02", X"14", X"40", X"00", X"69", 
  X"00", X"00", X"00", X"00", X"8c", X"a7", X"00", X"00", 
  X"2c", X"e2", X"00", X"02", X"14", X"40", X"00", X"63", 
  X"00", X"a0", X"10", X"21", X"24", X"02", X"00", X"04", 
  X"10", X"62", X"00", X"64", X"00", X"00", X"00", X"00", 
  X"10", X"e2", X"00", X"5e", X"00", X"a0", X"10", X"21", 
  X"24", X"02", X"00", X"02", X"10", X"e2", X"00", X"5d", 
  X"00", X"00", X"00", X"00", X"10", X"62", X"00", X"59", 
  X"00", X"a0", X"10", X"21", X"8c", X"83", X"00", X"08", 
  X"8c", X"ac", X"00", X"08", X"8c", X"8b", X"00", X"10", 
  X"8c", X"88", X"00", X"14", X"00", X"6c", X"38", X"23", 
  X"00", X"07", X"17", X"c3", X"00", X"47", X"38", X"26", 
  X"00", X"e2", X"10", X"23", X"28", X"42", X"00", X"40", 
  X"8c", X"aa", X"00", X"10", X"14", X"40", X"00", X"5a", 
  X"8c", X"a9", X"00", X"14", X"01", X"83", X"10", X"2a", 
  X"10", X"40", X"00", X"80", X"00", X"00", X"00", X"00", 
  X"00", X"60", X"60", X"21", X"00", X"00", X"50", X"21", 
  X"00", X"00", X"48", X"21", X"8c", X"82", X"00", X"04", 
  X"8c", X"a3", X"00", X"04", X"10", X"43", X"00", X"71", 
  X"01", X"09", X"18", X"21", X"10", X"40", X"00", X"6b", 
  X"01", X"09", X"18", X"23", X"01", X"28", X"18", X"23", 
  X"01", X"23", X"48", X"2b", X"01", X"4b", X"28", X"23", 
  X"00", X"a9", X"28", X"23", X"18", X"a0", X"00", X"74", 
  X"00", X"00", X"00", X"00", X"ac", X"c0", X"00", X"04", 
  X"ac", X"cc", X"00", X"08", X"ac", X"c5", X"00", X"10", 
  X"ac", X"c3", X"00", X"14", X"24", X"67", X"ff", X"ff", 
  X"00", X"e3", X"20", X"2b", X"24", X"a2", X"ff", X"ff", 
  X"00", X"82", X"10", X"21", X"3c", X"04", X"10", X"00", 
  X"00", X"44", X"40", X"2b", X"11", X"00", X"00", X"1d", 
  X"24", X"84", X"ff", X"ff", X"10", X"44", X"00", X"74", 
  X"00", X"00", X"00", X"00", X"8c", X"c7", X"00", X"08", 
  X"3c", X"04", X"10", X"00", X"00", X"a0", X"40", X"21", 
  X"24", X"e7", X"ff", X"ff", X"0b", X"f0", X"02", X"ef", 
  X"24", X"8d", X"ff", X"ff", X"11", X"2d", X"00", X"4b", 
  X"2d", X"4a", X"ff", X"ff", X"00", X"03", X"17", X"c2", 
  X"00", X"03", X"60", X"40", X"00", X"08", X"28", X"40", 
  X"00", X"45", X"28", X"25", X"25", X"8a", X"ff", X"ff", 
  X"24", X"a2", X"ff", X"ff", X"01", X"4c", X"48", X"2b", 
  X"01", X"22", X"48", X"21", X"01", X"24", X"10", X"2b", 
  X"00", X"e0", X"58", X"21", X"01", X"80", X"18", X"21", 
  X"00", X"a0", X"40", X"21", X"14", X"40", X"ff", X"f1", 
  X"24", X"e7", X"ff", X"ff", X"ac", X"c5", X"00", X"10", 
  X"ac", X"cc", X"00", X"14", X"ac", X"cb", X"00", X"08", 
  X"01", X"80", X"18", X"21", X"3c", X"02", X"20", X"00", 
  X"24", X"04", X"00", X"03", X"00", X"a2", X"10", X"2b", 
  X"14", X"40", X"00", X"0c", X"ac", X"c4", X"00", X"00", 
  X"8c", X"c4", X"00", X"08", X"00", X"05", X"3f", X"c0", 
  X"00", X"03", X"10", X"42", X"00", X"e2", X"10", X"25", 
  X"30", X"63", X"00", X"01", X"00", X"05", X"28", X"42", 
  X"00", X"43", X"10", X"25", X"24", X"84", X"00", X"01", 
  X"ac", X"c5", X"00", X"10", X"ac", X"c2", X"00", X"14", 
  X"ac", X"c4", X"00", X"08", X"03", X"e0", X"00", X"08", 
  X"00", X"c0", X"10", X"21", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"80", X"10", X"21", X"14", X"e3", X"ff", X"fb", 
  X"00", X"80", X"10", X"21", X"8c", X"84", X"00", X"04", 
  X"8c", X"a3", X"00", X"04", X"10", X"83", X"ff", X"f7", 
  X"00", X"00", X"00", X"00", X"3c", X"02", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"42", X"08", X"b0", 
  X"01", X"83", X"10", X"2a", X"10", X"40", X"00", X"0b", 
  X"00", X"6c", X"10", X"2a", X"00", X"0a", X"17", X"c0", 
  X"00", X"09", X"38", X"42", X"00", X"47", X"38", X"25", 
  X"31", X"29", X"00", X"01", X"25", X"8c", X"00", X"01", 
  X"00", X"0a", X"50", X"42", X"15", X"83", X"ff", X"f9", 
  X"00", X"e9", X"48", X"25", X"00", X"60", X"60", X"21", 
  X"00", X"6c", X"10", X"2a", X"10", X"40", X"00", X"31", 
  X"00", X"00", X"00", X"00", X"00", X"0b", X"17", X"c0", 
  X"00", X"08", X"38", X"42", X"00", X"47", X"38", X"25", 
  X"31", X"08", X"00", X"01", X"24", X"63", X"00", X"01", 
  X"00", X"0b", X"58", X"42", X"14", X"6c", X"ff", X"f9", 
  X"00", X"e8", X"40", X"25", X"0b", X"f0", X"02", X"ce", 
  X"8c", X"82", X"00", X"04", X"15", X"40", X"ff", X"b6", 
  X"00", X"03", X"17", X"c2", X"0b", X"f0", X"02", X"fe", 
  X"ac", X"c5", X"00", X"10", X"01", X"03", X"40", X"2b", 
  X"01", X"6a", X"28", X"23", X"0b", X"f0", X"02", X"d7", 
  X"00", X"a8", X"28", X"23", X"00", X"68", X"28", X"2b", 
  X"01", X"6a", X"50", X"21", X"00", X"aa", X"28", X"21", 
  X"ac", X"c2", X"00", X"04", X"ac", X"cc", X"00", X"08", 
  X"ac", X"c5", X"00", X"10", X"0b", X"f0", X"03", X"01", 
  X"ac", X"c3", X"00", X"14", X"00", X"00", X"58", X"21", 
  X"0b", X"f0", X"02", X"cd", X"00", X"00", X"40", X"21", 
  X"14", X"a0", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"14", X"60", X"ff", X"8a", X"00", X"00", X"00", X"00", 
  X"00", X"03", X"18", X"23", X"00", X"03", X"10", X"2b", 
  X"00", X"05", X"28", X"23", X"00", X"a2", X"28", X"23", 
  X"24", X"02", X"00", X"01", X"ac", X"c2", X"00", X"04", 
  X"ac", X"cc", X"00", X"08", X"ac", X"c5", X"00", X"10", 
  X"0b", X"f0", X"02", X"dd", X"ac", X"c3", X"00", X"14", 
  X"2c", X"e7", X"ff", X"ff", X"14", X"e0", X"ff", X"8b", 
  X"3c", X"02", X"20", X"00", X"0b", X"f0", X"03", X"03", 
  X"24", X"04", X"00", X"03", X"0b", X"f0", X"02", X"cd", 
  X"00", X"60", X"60", X"21", X"27", X"bd", X"ff", X"a0", 
  X"af", X"a5", X"00", X"64", X"af", X"a4", X"00", X"60", 
  X"27", X"a5", X"00", X"40", X"27", X"a4", X"00", X"60", 
  X"af", X"bf", X"00", X"5c", X"af", X"a7", X"00", X"6c", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"68", 
  X"27", X"a4", X"00", X"68", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"40", 
  X"27", X"a5", X"00", X"28", X"0f", X"f0", X"02", X"a9", 
  X"27", X"a6", X"00", X"10", X"0f", X"f0", X"01", X"c9", 
  X"00", X"40", X"20", X"21", X"8f", X"bf", X"00", X"5c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"60", 
  X"27", X"bd", X"ff", X"a0", X"af", X"a5", X"00", X"64", 
  X"af", X"a4", X"00", X"60", X"27", X"a5", X"00", X"40", 
  X"27", X"a4", X"00", X"60", X"af", X"bf", X"00", X"5c", 
  X"af", X"a7", X"00", X"6c", X"0f", X"f0", X"02", X"25", 
  X"af", X"a6", X"00", X"68", X"27", X"a4", X"00", X"68", 
  X"0f", X"f0", X"02", X"25", X"27", X"a5", X"00", X"28", 
  X"8f", X"a2", X"00", X"2c", X"27", X"a4", X"00", X"40", 
  X"27", X"a5", X"00", X"28", X"27", X"a6", X"00", X"10", 
  X"38", X"42", X"00", X"01", X"0f", X"f0", X"02", X"a9", 
  X"af", X"a2", X"00", X"2c", X"0f", X"f0", X"01", X"c9", 
  X"00", X"40", X"20", X"21", X"8f", X"bf", X"00", X"5c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"60", 
  X"27", X"bd", X"ff", X"a0", X"af", X"a5", X"00", X"64", 
  X"af", X"a4", X"00", X"60", X"27", X"a5", X"00", X"40", 
  X"27", X"a4", X"00", X"60", X"af", X"bf", X"00", X"5c", 
  X"af", X"a7", X"00", X"6c", X"0f", X"f0", X"02", X"25", 
  X"af", X"a6", X"00", X"68", X"27", X"a4", X"00", X"68", 
  X"0f", X"f0", X"02", X"25", X"27", X"a5", X"00", X"28", 
  X"8f", X"a2", X"00", X"40", X"2c", X"43", X"00", X"02", 
  X"14", X"60", X"00", X"72", X"8f", X"a3", X"00", X"28", 
  X"2c", X"64", X"00", X"02", X"14", X"80", X"00", X"7d", 
  X"24", X"04", X"00", X"04", X"10", X"44", X"00", X"6a", 
  X"00", X"00", X"00", X"00", X"10", X"64", X"00", X"76", 
  X"24", X"04", X"00", X"02", X"10", X"44", X"00", X"69", 
  X"00", X"00", X"00", X"00", X"10", X"64", X"00", X"75", 
  X"8f", X"a4", X"00", X"54", X"8f", X"a9", X"00", X"38", 
  X"8f", X"a8", X"00", X"50", X"8f", X"a5", X"00", X"3c", 
  X"01", X"24", X"00", X"19", X"00", X"00", X"10", X"10", 
  X"00", X"00", X"18", X"12", X"00", X"a8", X"00", X"19", 
  X"00", X"00", X"38", X"12", X"00", X"e3", X"50", X"21", 
  X"01", X"47", X"38", X"2b", X"00", X"00", X"30", X"10", 
  X"00", X"c2", X"30", X"21", X"00", X"e6", X"30", X"21", 
  X"00", X"a4", X"00", X"19", X"00", X"c2", X"38", X"2b", 
  X"00", X"00", X"28", X"12", X"00", X"00", X"20", X"10", 
  X"01", X"28", X"00", X"19", X"00", X"00", X"48", X"12", 
  X"10", X"e0", X"00", X"6a", X"00", X"00", X"40", X"10", 
  X"24", X"0b", X"00", X"01", X"01", X"44", X"18", X"21", 
  X"00", X"c9", X"38", X"21", X"00", X"64", X"10", X"2b", 
  X"8f", X"a9", X"00", X"48", X"8f", X"a4", X"00", X"30", 
  X"00", X"e6", X"30", X"2b", X"8f", X"aa", X"00", X"44", 
  X"01", X"24", X"48", X"21", X"8f", X"a4", X"00", X"2c", 
  X"00", X"c8", X"40", X"21", X"00", X"e2", X"10", X"21", 
  X"00", X"47", X"38", X"2b", X"01", X"0b", X"40", X"21", 
  X"00", X"e8", X"40", X"21", X"01", X"44", X"50", X"26", 
  X"3c", X"06", X"20", X"00", X"00", X"0a", X"50", X"2b", 
  X"25", X"27", X"00", X"04", X"01", X"06", X"30", X"2b", 
  X"00", X"a0", X"20", X"21", X"af", X"aa", X"00", X"14", 
  X"af", X"a7", X"00", X"18", X"25", X"25", X"00", X"05", 
  X"3c", X"0f", X"80", X"00", X"14", X"c0", X"00", X"11", 
  X"3c", X"0d", X"20", X"00", X"00", X"08", X"3f", X"c0", 
  X"30", X"49", X"00", X"01", X"00", X"08", X"40", X"42", 
  X"00", X"02", X"10", X"42", X"01", X"0d", X"30", X"2b", 
  X"00", X"03", X"5f", X"c0", X"00", X"04", X"50", X"42", 
  X"00", X"03", X"60", X"42", X"11", X"20", X"00", X"03", 
  X"00", X"a0", X"70", X"21", X"01", X"8f", X"18", X"25", 
  X"01", X"6a", X"20", X"25", X"00", X"e2", X"10", X"25", 
  X"10", X"c0", X"ff", X"f2", X"24", X"a5", X"00", X"01", 
  X"af", X"ae", X"00", X"18", X"3c", X"05", X"10", X"00", 
  X"01", X"05", X"28", X"2b", X"10", X"a0", X"00", X"13", 
  X"8f", X"a5", X"00", X"18", X"3c", X"0c", X"10", X"00", 
  X"24", X"a5", X"ff", X"ff", X"00", X"02", X"37", X"c2", 
  X"00", X"08", X"40", X"40", X"00", X"02", X"10", X"40", 
  X"00", X"c8", X"40", X"25", X"28", X"6a", X"00", X"00", 
  X"00", X"04", X"3f", X"c2", X"34", X"49", X"00", X"01", 
  X"00", X"03", X"18", X"40", X"01", X"0c", X"30", X"2b", 
  X"00", X"a0", X"58", X"21", X"01", X"2a", X"10", X"0b", 
  X"00", X"e3", X"18", X"25", X"00", X"04", X"20", X"40", 
  X"14", X"c0", X"ff", X"f2", X"24", X"a5", X"ff", X"ff", 
  X"af", X"ab", X"00", X"18", X"30", X"46", X"00", X"ff", 
  X"24", X"05", X"00", X"80", X"10", X"c5", X"00", X"2e", 
  X"30", X"45", X"01", X"00", X"af", X"a2", X"00", X"24", 
  X"27", X"a4", X"00", X"10", X"24", X"02", X"00", X"03", 
  X"af", X"a8", X"00", X"20", X"0f", X"f0", X"01", X"c9", 
  X"af", X"a2", X"00", X"10", X"8f", X"bf", X"00", X"5c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"60", 
  X"24", X"02", X"00", X"02", X"10", X"62", X"00", X"20", 
  X"3c", X"04", X"00", X"00", X"8f", X"a3", X"00", X"44", 
  X"8f", X"a2", X"00", X"2c", X"27", X"a4", X"00", X"40", 
  X"00", X"62", X"10", X"26", X"00", X"02", X"10", X"2b", 
  X"af", X"a2", X"00", X"44", X"0f", X"f0", X"01", X"c9", 
  X"00", X"00", X"00", X"00", X"8f", X"bf", X"00", X"5c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"60", 
  X"24", X"03", X"00", X"02", X"10", X"43", X"00", X"12", 
  X"3c", X"04", X"00", X"00", X"8f", X"a2", X"00", X"2c", 
  X"8f", X"a3", X"00", X"44", X"27", X"a4", X"00", X"28", 
  X"00", X"62", X"10", X"26", X"00", X"02", X"10", X"2b", 
  X"0f", X"f0", X"01", X"c9", X"af", X"a2", X"00", X"2c", 
  X"8f", X"bf", X"00", X"5c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"60", X"14", X"c2", X"ff", X"97", 
  X"00", X"00", X"58", X"21", X"01", X"43", X"10", X"2b", 
  X"14", X"40", X"ff", X"93", X"01", X"44", X"18", X"21", 
  X"0b", X"f0", X"03", X"c0", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"04", X"15", X"24", X"84", X"08", X"b0", 
  X"14", X"a0", X"00", X"03", X"00", X"64", X"18", X"25", 
  X"10", X"60", X"ff", X"d0", X"00", X"00", X"00", X"00", 
  X"24", X"43", X"00", X"80", X"00", X"62", X"10", X"2b", 
  X"00", X"48", X"40", X"21", X"0b", X"f0", X"04", X"03", 
  X"00", X"60", X"10", X"21", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"8f", X"a2", X"00", X"28", 
  X"2c", X"43", X"00", X"02", X"14", X"60", X"00", X"56", 
  X"8f", X"a3", X"00", X"10", X"2c", X"64", X"00", X"02", 
  X"14", X"80", X"00", X"58", X"8f", X"a6", X"00", X"2c", 
  X"8f", X"a5", X"00", X"14", X"24", X"04", X"00", X"04", 
  X"00", X"c5", X"28", X"26", X"10", X"44", X"00", X"40", 
  X"af", X"a5", X"00", X"2c", X"24", X"05", X"00", X"02", 
  X"10", X"45", X"00", X"3d", X"00", X"00", X"00", X"00", 
  X"10", X"64", X"00", X"56", X"00", X"00", X"10", X"21", 
  X"10", X"65", X"00", X"63", X"8f", X"a2", X"00", X"18", 
  X"8f", X"a4", X"00", X"30", X"8f", X"a3", X"00", X"38", 
  X"8f", X"a7", X"00", X"20", X"00", X"82", X"20", X"23", 
  X"af", X"a4", X"00", X"30", X"00", X"67", X"40", X"2b", 
  X"8f", X"a2", X"00", X"3c", X"11", X"00", X"00", X"37", 
  X"8f", X"ad", X"00", X"24", X"00", X"02", X"2f", X"c2", 
  X"00", X"03", X"18", X"40", X"00", X"a3", X"18", X"25", 
  X"24", X"84", X"ff", X"ff", X"00", X"02", X"10", X"40", 
  X"af", X"a4", X"00", X"30", X"00", X"67", X"40", X"2b", 
  X"24", X"05", X"00", X"3d", X"3c", X"04", X"10", X"00", 
  X"00", X"00", X"30", X"21", X"00", X"00", X"60", X"21", 
  X"0b", X"f0", X"04", X"6f", X"00", X"00", X"58", X"21", 
  X"00", X"67", X"40", X"2b", X"00", X"04", X"57", X"c0", 
  X"00", X"06", X"48", X"42", X"15", X"00", X"00", X"0c", 
  X"24", X"a5", X"ff", X"ff", X"00", X"4d", X"40", X"23", 
  X"00", X"48", X"70", X"2b", X"00", X"67", X"78", X"23", 
  X"14", X"e3", X"00", X"03", X"00", X"4d", X"c0", X"2b", 
  X"17", X"00", X"00", X"05", X"00", X"00", X"00", X"00", 
  X"01", X"ee", X"18", X"23", X"01", X"00", X"10", X"21", 
  X"01", X"84", X"60", X"25", X"01", X"66", X"58", X"25", 
  X"00", X"02", X"37", X"c2", X"00", X"03", X"18", X"40", 
  X"00", X"c3", X"18", X"25", X"00", X"04", X"20", X"42", 
  X"01", X"49", X"30", X"25", X"14", X"a0", X"ff", X"ea", 
  X"00", X"02", X"10", X"40", X"31", X"65", X"00", X"ff", 
  X"24", X"04", X"00", X"80", X"10", X"a4", X"00", X"29", 
  X"31", X"64", X"01", X"00", X"27", X"a4", X"00", X"28", 
  X"af", X"ac", X"00", X"38", X"0f", X"f0", X"01", X"c9", 
  X"af", X"ab", X"00", X"3c", X"8f", X"bf", X"00", X"44", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"48", 
  X"10", X"43", X"00", X"17", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"01", X"c9", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"14", X"e3", X"ff", X"d1", 
  X"24", X"05", X"00", X"3d", X"00", X"4d", X"28", X"2b", 
  X"10", X"a0", X"ff", X"cd", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"04", X"62", X"00", X"02", X"2f", X"c2", 
  X"0f", X"f0", X"01", X"c9", X"27", X"a4", X"00", X"28", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"0f", X"f0", X"01", X"c9", 
  X"27", X"a4", X"00", X"10", X"8f", X"bf", X"00", X"44", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"48", 
  X"3c", X"04", X"00", X"00", X"0b", X"f0", X"04", X"92", 
  X"24", X"84", X"08", X"b0", X"00", X"00", X"18", X"21", 
  X"af", X"a3", X"00", X"3c", X"af", X"a2", X"00", X"38", 
  X"af", X"a0", X"00", X"30", X"0b", X"f0", X"04", X"92", 
  X"27", X"a4", X"00", X"28", X"14", X"80", X"00", X"03", 
  X"00", X"62", X"10", X"25", X"10", X"40", X"ff", X"d6", 
  X"27", X"a4", X"00", X"28", X"25", X"62", X"00", X"80", 
  X"00", X"4b", X"58", X"2b", X"01", X"6c", X"60", X"21", 
  X"0b", X"f0", X"04", X"89", X"00", X"40", X"58", X"21", 
  X"af", X"a4", X"00", X"28", X"0b", X"f0", X"04", X"92", 
  X"27", X"a4", X"00", X"10", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"02", X"60", X"27", X"a5", X"00", X"10", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"8f", X"a2", X"00", X"28", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"09", 
  X"8f", X"a2", X"00", X"10", X"2c", X"42", X"00", X"02", 
  X"14", X"40", X"00", X"06", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"02", X"60", X"27", X"a5", X"00", X"10", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"8f", X"bf", X"00", X"44", 
  X"24", X"02", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"8f", X"a2", X"00", X"28", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"09", 
  X"8f", X"a2", X"00", X"10", X"2c", X"42", X"00", X"02", 
  X"14", X"40", X"00", X"06", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"02", X"60", X"27", X"a5", X"00", X"10", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"8f", X"bf", X"00", X"44", 
  X"24", X"02", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"8f", X"a2", X"00", X"28", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"07", 
  X"24", X"02", X"ff", X"ff", X"8f", X"a2", X"00", X"10", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"06", 
  X"27", X"a4", X"00", X"28", X"0f", X"f0", X"02", X"60", 
  X"27", X"a5", X"00", X"10", X"8f", X"bf", X"00", X"44", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"48", 
  X"0b", X"f0", X"05", X"1d", X"24", X"02", X"ff", X"ff", 
  X"27", X"bd", X"ff", X"b8", X"af", X"a5", X"00", X"4c", 
  X"af", X"a4", X"00", X"48", X"27", X"a5", X"00", X"28", 
  X"27", X"a4", X"00", X"48", X"af", X"bf", X"00", X"44", 
  X"af", X"a7", X"00", X"54", X"0f", X"f0", X"02", X"25", 
  X"af", X"a6", X"00", X"50", X"27", X"a4", X"00", X"50", 
  X"0f", X"f0", X"02", X"25", X"27", X"a5", X"00", X"10", 
  X"8f", X"a2", X"00", X"28", X"2c", X"42", X"00", X"02", 
  X"14", X"40", X"00", X"07", X"24", X"02", X"ff", X"ff", 
  X"8f", X"a2", X"00", X"10", X"2c", X"42", X"00", X"02", 
  X"14", X"40", X"00", X"06", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"02", X"60", X"27", X"a5", X"00", X"10", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"0b", X"f0", X"05", X"38", 
  X"24", X"02", X"ff", X"ff", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"8f", X"a2", X"00", X"28", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"09", 
  X"8f", X"a2", X"00", X"10", X"2c", X"42", X"00", X"02", 
  X"14", X"40", X"00", X"06", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"02", X"60", X"27", X"a5", X"00", X"10", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"8f", X"bf", X"00", X"44", 
  X"24", X"02", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"27", X"bd", X"ff", X"b8", 
  X"af", X"a5", X"00", X"4c", X"af", X"a4", X"00", X"48", 
  X"27", X"a5", X"00", X"28", X"27", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"af", X"a7", X"00", X"54", 
  X"0f", X"f0", X"02", X"25", X"af", X"a6", X"00", X"50", 
  X"27", X"a4", X"00", X"50", X"0f", X"f0", X"02", X"25", 
  X"27", X"a5", X"00", X"10", X"8f", X"a2", X"00", X"28", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"09", 
  X"8f", X"a2", X"00", X"10", X"2c", X"42", X"00", X"02", 
  X"14", X"40", X"00", X"06", X"27", X"a4", X"00", X"28", 
  X"0f", X"f0", X"02", X"60", X"27", X"a5", X"00", X"10", 
  X"8f", X"bf", X"00", X"44", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"8f", X"bf", X"00", X"44", 
  X"24", X"02", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"27", X"bd", X"ff", X"d0", 
  X"00", X"04", X"17", X"c2", X"24", X"03", X"00", X"03", 
  X"af", X"bf", X"00", X"2c", X"af", X"a3", X"00", X"10", 
  X"14", X"80", X"00", X"08", X"af", X"a2", X"00", X"14", 
  X"24", X"02", X"00", X"02", X"af", X"a2", X"00", X"10", 
  X"0f", X"f0", X"01", X"c9", X"27", X"a4", X"00", X"10", 
  X"8f", X"bf", X"00", X"2c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"24", X"03", X"00", X"3c", 
  X"14", X"40", X"00", X"15", X"af", X"a3", X"00", X"18", 
  X"00", X"04", X"17", X"c3", X"af", X"a2", X"00", X"20", 
  X"af", X"a4", X"00", X"24", X"3c", X"03", X"10", X"00", 
  X"00", X"43", X"18", X"2b", X"10", X"60", X"ff", X"f2", 
  X"24", X"03", X"00", X"3b", X"3c", X"07", X"10", X"00", 
  X"00", X"04", X"2f", X"c2", X"00", X"02", X"10", X"40", 
  X"00", X"a2", X"10", X"25", X"00", X"47", X"28", X"2b", 
  X"00", X"60", X"30", X"21", X"00", X"04", X"20", X"40", 
  X"14", X"a0", X"ff", X"f9", X"24", X"63", X"ff", X"ff", 
  X"af", X"a2", X"00", X"20", X"af", X"a4", X"00", X"24", 
  X"0b", X"f0", X"05", X"7e", X"af", X"a6", X"00", X"18", 
  X"3c", X"02", X"80", X"00", X"10", X"82", X"00", X"06", 
  X"3c", X"03", X"80", X"00", X"00", X"04", X"20", X"23", 
  X"00", X"04", X"17", X"c3", X"af", X"a2", X"00", X"20", 
  X"0b", X"f0", X"05", X"89", X"af", X"a4", X"00", X"24", 
  X"0b", X"f0", X"05", X"80", X"24", X"02", X"ff", X"ff", 
  X"27", X"bd", X"ff", X"d0", X"af", X"a5", X"00", X"34", 
  X"af", X"a4", X"00", X"30", X"27", X"a5", X"00", X"10", 
  X"af", X"bf", X"00", X"2c", X"0f", X"f0", X"02", X"25", 
  X"27", X"a4", X"00", X"30", X"8f", X"a2", X"00", X"10", 
  X"2c", X"43", X"00", X"03", X"14", X"60", X"00", X"0e", 
  X"24", X"03", X"00", X"04", X"10", X"43", X"00", X"05", 
  X"8f", X"a2", X"00", X"18", X"04", X"40", X"00", X"0a", 
  X"28", X"43", X"00", X"1f", X"14", X"60", X"00", X"0c", 
  X"24", X"03", X"00", X"3c", X"8f", X"a2", X"00", X"14", 
  X"14", X"40", X"00", X"1a", X"8f", X"bf", X"00", X"2c", 
  X"3c", X"02", X"7f", X"ff", X"34", X"42", X"ff", X"ff", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"8f", X"bf", X"00", X"2c", X"00", X"00", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"8f", X"a4", X"00", X"20", X"00", X"62", X"10", X"23", 
  X"00", X"02", X"18", X"27", X"00", X"04", X"30", X"40", 
  X"00", X"66", X"30", X"04", X"8f", X"a3", X"00", X"24", 
  X"30", X"45", X"00", X"20", X"8f", X"bf", X"00", X"2c", 
  X"00", X"43", X"18", X"06", X"00", X"c3", X"18", X"25", 
  X"00", X"44", X"10", X"06", X"8f", X"a4", X"00", X"14", 
  X"00", X"45", X"18", X"0b", X"00", X"03", X"10", X"23", 
  X"00", X"64", X"10", X"0a", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"3c", X"02", X"80", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"27", X"bd", X"ff", X"d0", X"af", X"a5", X"00", X"34", 
  X"af", X"a4", X"00", X"30", X"27", X"a5", X"00", X"10", 
  X"af", X"bf", X"00", X"2c", X"0f", X"f0", X"02", X"25", 
  X"27", X"a4", X"00", X"30", X"8f", X"a2", X"00", X"14", 
  X"27", X"a4", X"00", X"10", X"2c", X"42", X"00", X"01", 
  X"0f", X"f0", X"01", X"c9", X"af", X"a2", X"00", X"14", 
  X"8f", X"bf", X"00", X"2c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"3c", X"03", X"80", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"27", X"bd", X"ff", X"d0", X"af", X"a4", X"00", X"10", 
  X"27", X"a4", X"00", X"10", X"af", X"bf", X"00", X"2c", 
  X"af", X"a5", X"00", X"14", X"af", X"a6", X"00", X"18", 
  X"af", X"a7", X"00", X"24", X"0f", X"f0", X"01", X"c9", 
  X"af", X"a0", X"00", X"20", X"8f", X"bf", X"00", X"2c", 
  X"00", X"60", X"10", X"21", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"27", X"bd", X"ff", X"b8", 
  X"27", X"a5", X"00", X"28", X"af", X"a4", X"00", X"48", 
  X"af", X"bf", X"00", X"44", X"0f", X"f0", X"02", X"25", 
  X"27", X"a4", X"00", X"48", X"8f", X"a5", X"00", X"28", 
  X"8f", X"a3", X"00", X"3c", X"8f", X"a2", X"00", X"38", 
  X"af", X"a5", X"00", X"10", X"8f", X"a5", X"00", X"2c", 
  X"00", X"03", X"20", X"82", X"00", X"02", X"17", X"80", 
  X"af", X"a5", X"00", X"14", X"8f", X"a5", X"00", X"30", 
  X"00", X"82", X"10", X"25", X"00", X"03", X"1f", X"80", 
  X"27", X"a4", X"00", X"10", X"af", X"a5", X"00", X"18", 
  X"af", X"a2", X"00", X"20", X"0f", X"f0", X"01", X"c9", 
  X"af", X"a3", X"00", X"24", X"8f", X"bf", X"00", X"44", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"48", 
  X"27", X"bd", X"ff", X"d0", X"8f", X"a3", X"00", X"44", 
  X"8f", X"a2", X"00", X"40", X"af", X"a4", X"00", X"10", 
  X"27", X"a4", X"00", X"10", X"af", X"bf", X"00", X"2c", 
  X"af", X"a5", X"00", X"14", X"af", X"a6", X"00", X"18", 
  X"af", X"a3", X"00", X"24", X"0f", X"f0", X"01", X"c9", 
  X"af", X"a2", X"00", X"20", X"8f", X"bf", X"00", X"2c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"27", X"bd", X"ff", X"b8", X"af", X"a5", X"00", X"4c", 
  X"af", X"a4", X"00", X"48", X"27", X"a5", X"00", X"28", 
  X"af", X"bf", X"00", X"44", X"0f", X"f0", X"02", X"25", 
  X"27", X"a4", X"00", X"48", X"8f", X"a3", X"00", X"3c", 
  X"8f", X"a2", X"00", X"38", X"af", X"a0", X"00", X"20", 
  X"00", X"03", X"27", X"82", X"00", X"02", X"10", X"80", 
  X"00", X"44", X"10", X"25", X"7c", X"63", X"e8", X"00", 
  X"34", X"44", X"00", X"01", X"00", X"83", X"10", X"0b", 
  X"8f", X"a3", X"00", X"28", X"27", X"a4", X"00", X"10", 
  X"af", X"a2", X"00", X"24", X"af", X"a3", X"00", X"10", 
  X"8f", X"a3", X"00", X"2c", X"af", X"a3", X"00", X"14", 
  X"8f", X"a3", X"00", X"30", X"0f", X"f0", X"01", X"c9", 
  X"af", X"a3", X"00", X"18", X"8f", X"bf", X"00", X"44", 
  X"00", X"60", X"10", X"21", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"48", X"03", X"e0", X"00", X"08", 
  X"24", X"02", X"ff", X"ff", X"24", X"02", X"20", X"00", 
  X"ac", X"a2", X"00", X"04", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"10", X"21", X"03", X"e0", X"00", X"08", 
  X"24", X"02", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"10", X"21", X"03", X"e0", X"00", X"08", 
  X"24", X"02", X"ff", X"ff", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"10", X"21", X"3c", X"03", X"00", X"00", 
  X"8c", X"62", X"08", X"c8", X"10", X"40", X"00", X"08", 
  X"3c", X"05", X"00", X"02", X"00", X"44", X"20", X"21", 
  X"24", X"a5", X"00", X"01", X"00", X"85", X"28", X"2b", 
  X"10", X"a0", X"00", X"09", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"ac", X"64", X"08", X"c8", 
  X"3c", X"02", X"00", X"01", X"00", X"44", X"20", X"21", 
  X"24", X"a5", X"00", X"01", X"00", X"85", X"28", X"2b", 
  X"14", X"a0", X"ff", X"f9", X"ac", X"62", X"08", X"c8", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"90", X"a2", X"00", X"00", X"3c", X"03", X"20", X"00", 
  X"10", X"40", X"00", X"06", X"24", X"a5", X"00", X"01", 
  X"a0", X"62", X"00", X"00", X"24", X"a5", X"00", X"01", 
  X"90", X"a2", X"ff", X"ff", X"14", X"40", X"ff", X"fc", 
  X"00", X"00", X"00", X"00", X"24", X"03", X"00", X"0a", 
  X"3c", X"02", X"20", X"00", X"a0", X"43", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"00", X"01", 
  X"90", X"82", X"00", X"00", X"3c", X"03", X"20", X"00", 
  X"10", X"40", X"00", X"06", X"24", X"84", X"00", X"01", 
  X"a0", X"62", X"00", X"00", X"24", X"84", X"00", X"01", 
  X"90", X"82", X"ff", X"ff", X"14", X"40", X"ff", X"fc", 
  X"00", X"00", X"00", X"00", X"24", X"03", X"00", X"0a", 
  X"3c", X"02", X"20", X"00", X"a0", X"43", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"00", X"01", 
  X"00", X"a4", X"18", X"2b", X"10", X"60", X"00", X"06", 
  X"00", X"80", X"10", X"21", X"00", X"45", X"10", X"23", 
  X"00", X"a2", X"18", X"2b", X"14", X"60", X"ff", X"fe", 
  X"00", X"45", X"10", X"23", X"00", X"45", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"00", X"a4", X"10", X"2b", X"10", X"40", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"10", X"21", 
  X"00", X"85", X"20", X"23", X"00", X"a4", X"18", X"2b", 
  X"14", X"60", X"ff", X"fd", X"24", X"42", X"00", X"01", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"27", X"bd", X"ff", X"e0", X"3c", X"02", X"00", X"00", 
  X"af", X"a6", X"00", X"28", X"00", X"80", X"30", X"21", 
  X"8c", X"44", X"08", X"9c", X"af", X"a7", X"00", X"2c", 
  X"af", X"a5", X"00", X"24", X"8c", X"85", X"00", X"08", 
  X"27", X"a7", X"00", X"24", X"af", X"bf", X"00", X"1c", 
  X"0f", X"f0", X"06", X"e3", X"af", X"a7", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"27", X"bd", X"ff", X"e0", 
  X"af", X"a6", X"00", X"28", X"af", X"a7", X"00", X"2c", 
  X"00", X"a0", X"30", X"21", X"8c", X"85", X"00", X"08", 
  X"27", X"a7", X"00", X"28", X"af", X"bf", X"00", X"1c", 
  X"0f", X"f0", X"06", X"e3", X"af", X"a7", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"8c", X"c2", X"00", X"08", 
  X"27", X"bd", X"ff", X"c8", X"af", X"b0", X"00", X"14", 
  X"af", X"bf", X"00", X"34", X"af", X"b7", X"00", X"30", 
  X"af", X"b6", X"00", X"2c", X"af", X"b5", X"00", X"28", 
  X"af", X"b4", X"00", X"24", X"af", X"b3", X"00", X"20", 
  X"af", X"b2", X"00", X"1c", X"af", X"b1", X"00", X"18", 
  X"10", X"40", X"00", X"26", X"00", X"c0", X"80", X"21", 
  X"8c", X"a2", X"00", X"60", X"30", X"42", X"20", X"00", 
  X"10", X"40", X"00", X"1c", X"00", X"a0", X"98", X"21", 
  X"8c", X"d1", X"00", X"00", X"00", X"80", X"a8", X"21", 
  X"24", X"16", X"ff", X"ff", X"8e", X"02", X"00", X"08", 
  X"10", X"40", X"00", X"1b", X"00", X"00", X"90", X"21", 
  X"8e", X"34", X"00", X"04", X"8e", X"37", X"00", X"00", 
  X"00", X"14", X"a0", X"82", X"02", X"54", X"10", X"2a", 
  X"10", X"40", X"00", X"0a", X"00", X"12", X"10", X"80", 
  X"02", X"e2", X"10", X"21", X"8c", X"45", X"00", X"00", 
  X"02", X"a0", X"20", X"21", X"0f", X"f0", X"0c", X"32", 
  X"02", X"60", X"30", X"21", X"10", X"56", X"00", X"0d", 
  X"26", X"52", X"00", X"01", X"0b", X"f0", X"06", X"c0", 
  X"02", X"54", X"10", X"2a", X"8e", X"02", X"00", X"08", 
  X"00", X"14", X"a0", X"80", X"26", X"31", X"00", X"08", 
  X"00", X"54", X"a0", X"23", X"0b", X"f0", X"06", X"b9", 
  X"ae", X"14", X"00", X"08", X"0f", X"f0", X"0d", X"8d", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"06", X"d7", 
  X"ae", X"00", X"00", X"08", X"24", X"02", X"ff", X"ff", 
  X"ae", X"00", X"00", X"08", X"8f", X"bf", X"00", X"34", 
  X"8f", X"b7", X"00", X"30", X"8f", X"b6", X"00", X"2c", 
  X"8f", X"b5", X"00", X"28", X"8f", X"b4", X"00", X"24", 
  X"8f", X"b3", X"00", X"20", X"8f", X"b2", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"ae", X"00", X"00", X"04", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"27", X"bd", X"ff", X"38", 
  X"af", X"be", X"00", X"c0", X"af", X"b2", X"00", X"a8", 
  X"af", X"b1", X"00", X"a4", X"af", X"bf", X"00", X"c4", 
  X"af", X"b7", X"00", X"bc", X"af", X"b6", X"00", X"b8", 
  X"af", X"b5", X"00", X"b4", X"af", X"b4", X"00", X"b0", 
  X"af", X"b3", X"00", X"ac", X"af", X"b0", X"00", X"a0", 
  X"00", X"80", X"90", X"21", X"00", X"a0", X"88", X"21", 
  X"af", X"a6", X"00", X"d0", X"10", X"80", X"00", X"06", 
  X"00", X"e0", X"f0", X"21", X"8c", X"82", X"00", X"38", 
  X"54", X"40", X"00", X"04", X"86", X"22", X"00", X"0c", 
  X"0f", X"f0", X"0b", X"91", X"00", X"00", X"00", X"00", 
  X"86", X"22", X"00", X"0c", X"30", X"43", X"20", X"00", 
  X"54", X"60", X"00", X"08", X"96", X"22", X"00", X"0c", 
  X"8e", X"23", X"00", X"60", X"34", X"42", X"20", X"00", 
  X"a6", X"22", X"00", X"0c", X"24", X"02", X"df", X"ff", 
  X"00", X"62", X"10", X"24", X"ae", X"22", X"00", X"60", 
  X"96", X"22", X"00", X"0c", X"30", X"42", X"00", X"08", 
  X"10", X"40", X"00", X"0b", X"02", X"40", X"20", X"21", 
  X"8e", X"22", X"00", X"10", X"10", X"40", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"96", X"23", X"00", X"0c", 
  X"24", X"02", X"00", X"0a", X"30", X"63", X"00", X"1a", 
  X"54", X"62", X"00", X"12", X"27", X"a2", X"00", X"10", 
  X"0b", X"f0", X"07", X"16", X"86", X"22", X"00", X"0e", 
  X"0f", X"f0", X"0a", X"69", X"02", X"20", X"28", X"21", 
  X"50", X"40", X"ff", X"f7", X"96", X"23", X"00", X"0c", 
  X"0b", X"f0", X"0a", X"25", X"24", X"02", X"ff", X"ff", 
  X"04", X"42", X"00", X"08", X"27", X"a2", X"00", X"10", 
  X"8f", X"a6", X"00", X"d0", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"0a", X"39", 
  X"03", X"c0", X"38", X"21", X"0b", X"f0", X"0a", X"26", 
  X"8f", X"bf", X"00", X"c4", X"af", X"a2", X"00", X"78", 
  X"af", X"a0", X"00", X"80", X"af", X"a0", X"00", X"7c", 
  X"00", X"40", X"48", X"21", X"af", X"a0", X"00", X"90", 
  X"af", X"a0", X"00", X"8c", X"8f", X"b0", X"00", X"d0", 
  X"24", X"03", X"00", X"25", X"92", X"02", X"00", X"00", 
  X"14", X"40", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"8f", X"a3", X"00", X"d0", X"02", X"03", X"a8", X"23", 
  X"56", X"a0", X"00", X"07", X"8f", X"a2", X"00", X"80", 
  X"0b", X"f0", X"07", X"49", X"92", X"02", X"00", X"00", 
  X"50", X"43", X"ff", X"fa", X"8f", X"a3", X"00", X"d0", 
  X"0b", X"f0", X"07", X"27", X"26", X"10", X"00", X"01", 
  X"8f", X"a4", X"00", X"d0", X"ad", X"35", X"00", X"04", 
  X"00", X"55", X"10", X"21", X"af", X"a2", X"00", X"80", 
  X"8f", X"a2", X"00", X"7c", X"ad", X"24", X"00", X"00", 
  X"24", X"42", X"00", X"01", X"af", X"a2", X"00", X"7c", 
  X"28", X"42", X"00", X"08", X"14", X"40", X"00", X"07", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"02", X"dc", 
  X"27", X"a9", X"00", X"10", X"8f", X"a5", X"00", X"8c", 
  X"00", X"b5", X"28", X"21", X"af", X"a5", X"00", X"8c", 
  X"92", X"02", X"00", X"00", X"10", X"40", X"02", X"cf", 
  X"26", X"03", X"00", X"01", X"a3", X"a0", X"00", X"86", 
  X"00", X"00", X"10", X"21", X"24", X"13", X"ff", X"ff", 
  X"af", X"a0", X"00", X"88", X"00", X"00", X"a0", X"21", 
  X"24", X"08", X"00", X"58", X"24", X"0a", X"00", X"2e", 
  X"24", X"06", X"00", X"2a", X"24", X"07", X"00", X"0a", 
  X"24", X"17", X"00", X"71", X"24", X"16", X"00", X"68", 
  X"24", X"15", X"00", X"69", X"24", X"0c", X"00", X"6c", 
  X"24", X"10", X"00", X"30", X"24", X"0e", X"00", X"2b", 
  X"24", X"0f", X"00", X"2d", X"24", X"0d", X"00", X"20", 
  X"24", X"18", X"00", X"23", X"24", X"64", X"00", X"01", 
  X"90", X"63", X"00", X"00", X"af", X"a4", X"00", X"d0", 
  X"10", X"68", X"00", X"5e", X"28", X"64", X"00", X"59", 
  X"10", X"80", X"00", X"2a", X"24", X"05", X"00", X"6e", 
  X"10", X"6a", X"00", X"66", X"8f", X"a5", X"00", X"d0", 
  X"28", X"64", X"00", X"2f", X"10", X"80", X"00", X"14", 
  X"28", X"64", X"00", X"3a", X"10", X"66", X"00", X"59", 
  X"28", X"64", X"00", X"2b", X"10", X"80", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"50", X"6d", X"00", X"04", 
  X"01", X"a2", X"10", X"0a", X"54", X"78", X"01", X"82", 
  X"a3", X"a2", X"00", X"86", X"36", X"94", X"00", X"01", 
  X"0b", X"f0", X"07", X"5d", X"8f", X"a3", X"00", X"d0", 
  X"14", X"6e", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"07", X"72", X"24", X"02", X"00", X"2b", 
  X"50", X"6f", X"ff", X"f9", X"36", X"94", X"00", X"04", 
  X"0b", X"f0", X"08", X"f2", X"a3", X"a2", X"00", X"86", 
  X"10", X"80", X"00", X"08", X"24", X"04", X"00", X"4f", 
  X"28", X"64", X"00", X"31", X"50", X"80", X"00", X"64", 
  X"af", X"a0", X"00", X"88", X"54", X"70", X"01", X"70", 
  X"a3", X"a2", X"00", X"86", X"0b", X"f0", X"07", X"72", 
  X"36", X"94", X"00", X"80", X"10", X"64", X"00", X"ad", 
  X"24", X"04", X"00", X"55", X"10", X"64", X"00", X"d6", 
  X"24", X"04", X"00", X"44", X"14", X"64", X"01", X"68", 
  X"a3", X"a2", X"00", X"86", X"0b", X"f0", X"08", X"00", 
  X"36", X"94", X"00", X"10", X"10", X"65", X"00", X"8f", 
  X"28", X"64", X"00", X"6f", X"10", X"80", X"00", X"12", 
  X"00", X"00", X"00", X"00", X"10", X"76", X"00", X"60", 
  X"28", X"64", X"00", X"69", X"10", X"80", X"00", X"08", 
  X"24", X"04", X"00", X"63", X"50", X"64", X"00", X"66", 
  X"8f", X"c2", X"00", X"00", X"24", X"04", X"00", X"64", 
  X"10", X"64", X"00", X"67", X"a3", X"a2", X"00", X"86", 
  X"0b", X"f0", X"08", X"f2", X"00", X"00", X"00", X"00", 
  X"50", X"75", X"00", X"63", X"a3", X"a2", X"00", X"86", 
  X"10", X"6c", X"00", X"55", X"8f", X"a4", X"00", X"d0", 
  X"0b", X"f0", X"08", X"f2", X"a3", X"a2", X"00", X"86", 
  X"10", X"77", X"00", X"57", X"28", X"64", X"00", X"72", 
  X"10", X"80", X"00", X"12", X"24", X"04", X"00", X"75", 
  X"24", X"04", X"00", X"6f", X"10", X"64", X"00", X"8c", 
  X"24", X"04", X"00", X"70", X"14", X"64", X"01", X"47", 
  X"00", X"00", X"b0", X"21", X"24", X"02", X"00", X"30", 
  X"a3", X"a2", X"00", X"84", X"24", X"02", X"00", X"78", 
  X"a3", X"a2", X"00", X"85", X"3c", X"02", X"bf", X"c0", 
  X"24", X"42", X"5c", X"e4", X"8f", X"d5", X"00", X"00", 
  X"af", X"a2", X"00", X"90", X"36", X"94", X"00", X"02", 
  X"27", X"de", X"00", X"04", X"0b", X"f0", X"08", X"97", 
  X"24", X"02", X"00", X"02", X"10", X"64", X"00", X"a7", 
  X"24", X"04", X"00", X"78", X"10", X"64", X"00", X"bb", 
  X"24", X"04", X"00", X"73", X"54", X"64", X"01", X"36", 
  X"a3", X"a2", X"00", X"86", X"0b", X"f0", X"08", X"4a", 
  X"8f", X"d0", X"00", X"00", X"a3", X"a2", X"00", X"86", 
  X"3c", X"02", X"bf", X"c0", X"0b", X"f0", X"08", X"78", 
  X"24", X"42", X"5c", X"d0", X"8f", X"c3", X"00", X"00", 
  X"27", X"de", X"00", X"04", X"04", X"61", X"ff", X"ac", 
  X"af", X"a3", X"00", X"88", X"00", X"03", X"18", X"23", 
  X"af", X"a3", X"00", X"88", X"0b", X"f0", X"07", X"72", 
  X"36", X"94", X"00", X"04", X"90", X"a3", X"00", X"00", 
  X"10", X"66", X"00", X"03", X"24", X"a4", X"00", X"01", 
  X"0b", X"f0", X"07", X"d7", X"00", X"00", X"28", X"21", 
  X"8f", X"d3", X"00", X"00", X"27", X"c3", X"00", X"04", 
  X"af", X"a4", X"00", X"d0", X"06", X"61", X"ff", X"9e", 
  X"00", X"60", X"f0", X"21", X"0b", X"f0", X"07", X"72", 
  X"24", X"13", X"ff", X"ff", X"24", X"6b", X"ff", X"d0", 
  X"2d", X"79", X"00", X"0a", X"53", X"20", X"00", X"06", 
  X"28", X"ab", X"00", X"00", X"70", X"a7", X"18", X"02", 
  X"24", X"84", X"00", X"01", X"00", X"6b", X"28", X"21", 
  X"0b", X"f0", X"07", X"d7", X"90", X"83", X"ff", X"ff", 
  X"24", X"13", X"ff", X"ff", X"00", X"ab", X"98", X"0a", 
  X"0b", X"f0", X"07", X"60", X"af", X"a4", X"00", X"d0", 
  X"8f", X"a4", X"00", X"88", X"24", X"63", X"ff", X"d0", 
  X"70", X"87", X"28", X"02", X"00", X"a3", X"20", X"21", 
  X"8f", X"a3", X"00", X"d0", X"af", X"a4", X"00", X"88", 
  X"24", X"64", X"00", X"01", X"90", X"83", X"ff", X"ff", 
  X"24", X"65", X"ff", X"d0", X"2c", X"a5", X"00", X"0a", 
  X"10", X"a0", X"ff", X"71", X"af", X"a4", X"00", X"d0", 
  X"0b", X"f0", X"07", X"e5", X"8f", X"a4", X"00", X"88", 
  X"0b", X"f0", X"07", X"72", X"36", X"94", X"00", X"40", 
  X"90", X"83", X"00", X"00", X"54", X"6c", X"ff", X"7c", 
  X"36", X"94", X"00", X"10", X"24", X"84", X"00", X"01", 
  X"0b", X"f0", X"07", X"fa", X"af", X"a4", X"00", X"d0", 
  X"0b", X"f0", X"07", X"72", X"36", X"94", X"00", X"20", 
  X"a3", X"a0", X"00", X"86", X"27", X"de", X"00", X"04", 
  X"0b", X"f0", X"08", X"f6", X"a3", X"a2", X"00", X"50", 
  X"32", X"82", X"00", X"20", X"10", X"40", X"00", X"08", 
  X"32", X"83", X"00", X"10", X"27", X"c8", X"00", X"07", 
  X"24", X"02", X"ff", X"f8", X"01", X"02", X"10", X"24", 
  X"24", X"5e", X"00", X"08", X"8c", X"56", X"00", X"00", 
  X"0b", X"f0", X"08", X"14", X"8c", X"55", X"00", X"04", 
  X"10", X"60", X"00", X"03", X"27", X"c2", X"00", X"04", 
  X"0b", X"f0", X"08", X"12", X"8f", X"d5", X"00", X"00", 
  X"32", X"83", X"00", X"40", X"10", X"60", X"00", X"02", 
  X"8f", X"d5", X"00", X"00", X"7c", X"15", X"ae", X"20", 
  X"00", X"15", X"b7", X"c3", X"00", X"40", X"f0", X"21", 
  X"06", X"c1", X"00", X"85", X"24", X"02", X"00", X"01", 
  X"00", X"15", X"a8", X"23", X"00", X"15", X"10", X"2b", 
  X"00", X"16", X"b0", X"23", X"02", X"c2", X"b0", X"23", 
  X"24", X"02", X"00", X"2d", X"0b", X"f0", X"08", X"99", 
  X"a3", X"a2", X"00", X"86", X"32", X"83", X"00", X"20", 
  X"a3", X"a2", X"00", X"86", X"10", X"60", X"00", X"06", 
  X"27", X"c2", X"00", X"04", X"8f", X"a5", X"00", X"8c", 
  X"8f", X"c3", X"00", X"00", X"00", X"05", X"27", X"c3", 
  X"0b", X"f0", X"08", X"30", X"ac", X"65", X"00", X"04", 
  X"32", X"83", X"00", X"10", X"14", X"60", X"00", X"07", 
  X"8f", X"c3", X"00", X"00", X"32", X"8a", X"00", X"40", 
  X"11", X"40", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"8f", X"a5", X"00", X"8c", X"0b", X"f0", X"08", X"31", 
  X"a4", X"65", X"00", X"00", X"8f", X"a4", X"00", X"8c", 
  X"ac", X"64", X"00", X"00", X"0b", X"f0", X"07", X"25", 
  X"00", X"40", X"f0", X"21", X"36", X"94", X"00", X"10", 
  X"32", X"82", X"00", X"20", X"10", X"40", X"00", X"08", 
  X"32", X"83", X"00", X"10", X"27", X"c8", X"00", X"07", 
  X"24", X"02", X"ff", X"f8", X"01", X"02", X"10", X"24", 
  X"24", X"5e", X"00", X"08", X"8c", X"56", X"00", X"00", 
  X"0b", X"f0", X"08", X"48", X"8c", X"55", X"00", X"04", 
  X"14", X"60", X"00", X"06", X"27", X"c2", X"00", X"04", 
  X"32", X"83", X"00", X"40", X"50", X"60", X"00", X"04", 
  X"8f", X"d5", X"00", X"00", X"0b", X"f0", X"08", X"46", 
  X"97", X"d5", X"00", X"02", X"8f", X"d5", X"00", X"00", 
  X"00", X"00", X"b0", X"21", X"00", X"40", X"f0", X"21", 
  X"0b", X"f0", X"08", X"97", X"00", X"00", X"10", X"21", 
  X"a3", X"a0", X"00", X"86", X"27", X"de", X"00", X"04", 
  X"06", X"60", X"00", X"0b", X"02", X"00", X"20", X"21", 
  X"00", X"00", X"28", X"21", X"02", X"60", X"30", X"21", 
  X"0f", X"f0", X"11", X"41", X"af", X"a9", X"00", X"98", 
  X"10", X"40", X"00", X"a7", X"8f", X"a9", X"00", X"98", 
  X"00", X"50", X"10", X"23", X"02", X"62", X"18", X"2a", 
  X"0b", X"f0", X"08", X"fa", X"00", X"43", X"98", X"0a", 
  X"0f", X"f0", X"14", X"dd", X"af", X"a9", X"00", X"98", 
  X"00", X"40", X"98", X"21", X"00", X"00", X"b0", X"21", 
  X"0b", X"f0", X"08", X"fb", X"8f", X"a9", X"00", X"98", 
  X"36", X"94", X"00", X"10", X"32", X"82", X"00", X"20", 
  X"10", X"40", X"00", X"08", X"32", X"83", X"00", X"10", 
  X"27", X"c8", X"00", X"07", X"24", X"02", X"ff", X"f8", 
  X"01", X"02", X"10", X"24", X"24", X"5e", X"00", X"08", 
  X"8c", X"56", X"00", X"00", X"0b", X"f0", X"08", X"73", 
  X"8c", X"55", X"00", X"04", X"14", X"60", X"00", X"06", 
  X"27", X"c2", X"00", X"04", X"32", X"83", X"00", X"40", 
  X"50", X"60", X"00", X"04", X"8f", X"d5", X"00", X"00", 
  X"0b", X"f0", X"08", X"71", X"97", X"d5", X"00", X"02", 
  X"8f", X"d5", X"00", X"00", X"00", X"00", X"b0", X"21", 
  X"00", X"40", X"f0", X"21", X"0b", X"f0", X"08", X"97", 
  X"24", X"02", X"00", X"01", X"a3", X"a2", X"00", X"86", 
  X"3c", X"02", X"bf", X"c0", X"24", X"42", X"5c", X"e4", 
  X"af", X"a2", X"00", X"90", X"32", X"82", X"00", X"20", 
  X"10", X"40", X"00", X"08", X"32", X"84", X"00", X"10", 
  X"27", X"c8", X"00", X"07", X"24", X"02", X"ff", X"f8", 
  X"01", X"02", X"10", X"24", X"24", X"5e", X"00", X"08", 
  X"8c", X"56", X"00", X"00", X"0b", X"f0", X"08", X"8d", 
  X"8c", X"55", X"00", X"04", X"14", X"80", X"00", X"06", 
  X"27", X"c2", X"00", X"04", X"32", X"84", X"00", X"40", 
  X"50", X"80", X"00", X"04", X"8f", X"d5", X"00", X"00", 
  X"0b", X"f0", X"08", X"8b", X"97", X"d5", X"00", X"02", 
  X"8f", X"d5", X"00", X"00", X"00", X"00", X"b0", X"21", 
  X"00", X"40", X"f0", X"21", X"32", X"84", X"00", X"01", 
  X"10", X"80", X"00", X"08", X"24", X"02", X"00", X"02", 
  X"02", X"d5", X"20", X"25", X"50", X"80", X"00", X"08", 
  X"a3", X"a0", X"00", X"86", X"24", X"04", X"00", X"30", 
  X"a3", X"a4", X"00", X"84", X"a3", X"a3", X"00", X"85", 
  X"36", X"94", X"00", X"02", X"0b", X"f0", X"08", X"9a", 
  X"a3", X"a0", X"00", X"86", X"24", X"02", X"00", X"01", 
  X"06", X"60", X"00", X"02", X"24", X"03", X"ff", X"7f", 
  X"02", X"83", X"a0", X"24", X"02", X"d5", X"18", X"25", 
  X"14", X"60", X"00", X"03", X"27", X"b7", X"00", X"78", 
  X"12", X"60", X"00", X"45", X"00", X"00", X"00", X"00", 
  X"24", X"03", X"00", X"01", X"10", X"43", X"00", X"16", 
  X"24", X"03", X"00", X"02", X"10", X"43", X"00", X"31", 
  X"02", X"e0", X"80", X"21", X"00", X"16", X"17", X"40", 
  X"32", X"a3", X"00", X"07", X"00", X"15", X"a8", X"c2", 
  X"00", X"16", X"b0", X"c2", X"00", X"55", X"a8", X"25", 
  X"26", X"10", X"ff", X"ff", X"24", X"63", X"00", X"30", 
  X"02", X"d5", X"10", X"25", X"14", X"40", X"ff", X"f7", 
  X"a2", X"03", X"00", X"00", X"32", X"82", X"00", X"01", 
  X"10", X"40", X"00", X"3b", X"02", X"00", X"20", X"21", 
  X"24", X"02", X"00", X"30", X"50", X"62", X"00", X"39", 
  X"02", X"60", X"b0", X"21", X"26", X"10", X"ff", X"ff", 
  X"0b", X"f0", X"08", X"ee", X"a0", X"82", X"ff", X"ff", 
  X"16", X"c0", X"00", X"07", X"02", X"e0", X"80", X"21", 
  X"2e", X"a2", X"00", X"0a", X"10", X"40", X"00", X"05", 
  X"02", X"c0", X"20", X"21", X"26", X"b5", X"00", X"30", 
  X"0b", X"f0", X"08", X"ed", X"a3", X"b5", X"00", X"77", 
  X"02", X"c0", X"20", X"21", X"02", X"a0", X"28", X"21", 
  X"24", X"07", X"00", X"0a", X"00", X"00", X"30", X"21", 
  X"0f", X"f0", X"06", X"74", X"af", X"a9", X"00", X"98", 
  X"24", X"63", X"00", X"30", X"26", X"10", X"ff", X"ff", 
  X"02", X"c0", X"20", X"21", X"02", X"a0", X"28", X"21", 
  X"a2", X"03", X"00", X"00", X"24", X"07", X"00", X"0a", 
  X"0f", X"f0", X"06", X"7e", X"00", X"00", X"30", X"21", 
  X"00", X"40", X"b0", X"21", X"00", X"62", X"10", X"25", 
  X"00", X"60", X"a8", X"21", X"14", X"40", X"ff", X"ee", 
  X"8f", X"a9", X"00", X"98", X"0b", X"f0", X"08", X"ef", 
  X"02", X"60", X"b0", X"21", X"8f", X"a5", X"00", X"90", 
  X"32", X"a2", X"00", X"0f", X"26", X"10", X"ff", X"ff", 
  X"00", X"a2", X"10", X"21", X"90", X"42", X"00", X"00", 
  X"00", X"15", X"a9", X"02", X"a2", X"02", X"00", X"00", 
  X"00", X"16", X"17", X"00", X"00", X"55", X"a8", X"25", 
  X"00", X"16", X"b1", X"02", X"02", X"d5", X"10", X"25", 
  X"14", X"40", X"ff", X"f5", X"8f", X"a5", X"00", X"90", 
  X"0b", X"f0", X"08", X"ef", X"02", X"60", X"b0", X"21", 
  X"14", X"40", X"00", X"07", X"02", X"e0", X"80", X"21", 
  X"32", X"82", X"00", X"01", X"50", X"40", X"00", X"05", 
  X"02", X"60", X"b0", X"21", X"24", X"02", X"00", X"30", 
  X"a3", X"a2", X"00", X"77", X"27", X"b0", X"00", X"77", 
  X"02", X"60", X"b0", X"21", X"0b", X"f0", X"08", X"fb", 
  X"02", X"f0", X"98", X"23", X"a3", X"a2", X"00", X"86", 
  X"10", X"60", X"01", X"27", X"8f", X"a2", X"00", X"80", 
  X"a3", X"a3", X"00", X"50", X"a3", X"a0", X"00", X"86", 
  X"24", X"13", X"00", X"01", X"00", X"00", X"b0", X"21", 
  X"0b", X"f0", X"08", X"fb", X"27", X"b0", X"00", X"50", 
  X"00", X"00", X"b0", X"21", X"02", X"76", X"a8", X"2a", 
  X"02", X"c0", X"10", X"21", X"02", X"75", X"10", X"0a", 
  X"00", X"40", X"a8", X"21", X"93", X"a2", X"00", X"86", 
  X"32", X"83", X"00", X"02", X"32", X"97", X"00", X"84", 
  X"00", X"02", X"10", X"2b", X"02", X"a2", X"a8", X"21", 
  X"af", X"a3", X"00", X"94", X"16", X"e0", X"00", X"33", 
  X"02", X"a3", X"a8", X"21", X"8f", X"a4", X"00", X"88", 
  X"00", X"95", X"18", X"23", X"18", X"60", X"00", X"2f", 
  X"24", X"07", X"00", X"10", X"28", X"65", X"00", X"11", 
  X"8f", X"a4", X"00", X"80", X"14", X"a0", X"00", X"19", 
  X"8f", X"a2", X"00", X"7c", X"3c", X"05", X"bf", X"c0", 
  X"24", X"42", X"00", X"01", X"24", X"a5", X"5c", X"50", 
  X"ad", X"25", X"00", X"00", X"24", X"84", X"00", X"10", 
  X"af", X"a2", X"00", X"7c", X"28", X"42", X"00", X"08", 
  X"ad", X"27", X"00", X"04", X"10", X"40", X"00", X"03", 
  X"af", X"a4", X"00", X"80", X"0b", X"f0", X"09", X"25", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"27", X"a6", X"00", X"78", 
  X"af", X"a3", X"00", X"98", X"0f", X"f0", X"06", X"a5", 
  X"af", X"a7", X"00", X"9c", X"8f", X"a3", X"00", X"98", 
  X"14", X"40", X"00", X"fd", X"8f", X"a7", X"00", X"9c", 
  X"27", X"a9", X"00", X"10", X"0b", X"f0", X"09", X"0b", 
  X"24", X"63", X"ff", X"f0", X"3c", X"05", X"bf", X"c0", 
  X"24", X"42", X"00", X"01", X"24", X"a5", X"5c", X"50", 
  X"ad", X"25", X"00", X"00", X"ad", X"23", X"00", X"04", 
  X"af", X"a2", X"00", X"7c", X"00", X"83", X"18", X"21", 
  X"28", X"42", X"00", X"08", X"10", X"40", X"00", X"03", 
  X"af", X"a3", X"00", X"80", X"0b", X"f0", X"09", X"39", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"00", X"e8", 
  X"27", X"a9", X"00", X"10", X"93", X"a2", X"00", X"86", 
  X"10", X"40", X"00", X"15", X"8f", X"a3", X"00", X"94", 
  X"27", X"a2", X"00", X"86", X"ad", X"22", X"00", X"00", 
  X"24", X"02", X"00", X"01", X"ad", X"22", X"00", X"04", 
  X"8f", X"a2", X"00", X"80", X"24", X"42", X"00", X"01", 
  X"af", X"a2", X"00", X"80", X"8f", X"a2", X"00", X"7c", 
  X"24", X"42", X"00", X"01", X"af", X"a2", X"00", X"7c", 
  X"28", X"42", X"00", X"08", X"14", X"40", X"00", X"07", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"00", X"d2", 
  X"27", X"a9", X"00", X"10", X"8f", X"a3", X"00", X"94", 
  X"10", X"60", X"00", X"15", X"24", X"02", X"00", X"80", 
  X"27", X"a2", X"00", X"84", X"ad", X"22", X"00", X"00", 
  X"24", X"02", X"00", X"02", X"ad", X"22", X"00", X"04", 
  X"8f", X"a2", X"00", X"80", X"24", X"42", X"00", X"02", 
  X"af", X"a2", X"00", X"80", X"8f", X"a2", X"00", X"7c", 
  X"24", X"42", X"00", X"01", X"af", X"a2", X"00", X"7c", 
  X"28", X"42", X"00", X"08", X"14", X"40", X"00", X"07", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"00", X"bc", 
  X"27", X"a9", X"00", X"10", X"24", X"02", X"00", X"80", 
  X"56", X"e2", X"00", X"32", X"02", X"d3", X"b0", X"23", 
  X"8f", X"a4", X"00", X"88", X"00", X"95", X"b8", X"23", 
  X"1a", X"e0", X"00", X"2d", X"24", X"07", X"00", X"10", 
  X"2a", X"e4", X"00", X"11", X"8f", X"a3", X"00", X"80", 
  X"14", X"80", X"00", X"17", X"8f", X"a2", X"00", X"7c", 
  X"24", X"42", X"00", X"01", X"3c", X"05", X"bf", X"c0", 
  X"24", X"a5", X"5c", X"40", X"24", X"63", X"00", X"10", 
  X"af", X"a2", X"00", X"7c", X"28", X"42", X"00", X"08", 
  X"ad", X"25", X"00", X"00", X"ad", X"27", X"00", X"04", 
  X"10", X"40", X"00", X"03", X"af", X"a3", X"00", X"80", 
  X"0b", X"f0", X"09", X"84", X"25", X"29", X"00", X"08", 
  X"02", X"40", X"20", X"21", X"02", X"20", X"28", X"21", 
  X"27", X"a6", X"00", X"78", X"0f", X"f0", X"06", X"a5", 
  X"af", X"a7", X"00", X"9c", X"14", X"40", X"00", X"9e", 
  X"8f", X"a7", X"00", X"9c", X"27", X"a9", X"00", X"10", 
  X"0b", X"f0", X"09", X"6c", X"26", X"f7", X"ff", X"f0", 
  X"24", X"42", X"00", X"01", X"3c", X"04", X"bf", X"c0", 
  X"24", X"84", X"5c", X"40", X"ad", X"37", X"00", X"04", 
  X"af", X"a2", X"00", X"7c", X"00", X"77", X"b8", X"21", 
  X"28", X"42", X"00", X"08", X"ad", X"24", X"00", X"00", 
  X"10", X"40", X"00", X"03", X"af", X"b7", X"00", X"80", 
  X"0b", X"f0", X"09", X"98", X"25", X"29", X"00", X"08", 
  X"02", X"40", X"20", X"21", X"02", X"20", X"28", X"21", 
  X"0f", X"f0", X"06", X"a5", X"27", X"a6", X"00", X"78", 
  X"14", X"40", X"00", X"89", X"27", X"a9", X"00", X"10", 
  X"02", X"d3", X"b0", X"23", X"1a", X"c0", X"00", X"2b", 
  X"24", X"17", X"00", X"10", X"2a", X"c4", X"00", X"11", 
  X"8f", X"a3", X"00", X"80", X"14", X"80", X"00", X"15", 
  X"8f", X"a2", X"00", X"7c", X"24", X"42", X"00", X"01", 
  X"3c", X"05", X"bf", X"c0", X"24", X"a5", X"5c", X"40", 
  X"24", X"63", X"00", X"10", X"af", X"a2", X"00", X"7c", 
  X"28", X"42", X"00", X"08", X"ad", X"25", X"00", X"00", 
  X"ad", X"37", X"00", X"04", X"10", X"40", X"00", X"03", 
  X"af", X"a3", X"00", X"80", X"0b", X"f0", X"09", X"b1", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"00", X"70", 
  X"27", X"a9", X"00", X"10", X"0b", X"f0", X"09", X"9b", 
  X"26", X"d6", X"ff", X"f0", X"24", X"42", X"00", X"01", 
  X"3c", X"04", X"bf", X"c0", X"24", X"84", X"5c", X"40", 
  X"ad", X"36", X"00", X"04", X"af", X"a2", X"00", X"7c", 
  X"00", X"76", X"b0", X"21", X"28", X"42", X"00", X"08", 
  X"ad", X"24", X"00", X"00", X"10", X"40", X"00", X"03", 
  X"af", X"b6", X"00", X"80", X"0b", X"f0", X"09", X"c5", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"00", X"5c", 
  X"27", X"a9", X"00", X"10", X"8f", X"a2", X"00", X"80", 
  X"ad", X"30", X"00", X"00", X"ad", X"33", X"00", X"04", 
  X"00", X"53", X"58", X"21", X"8f", X"a2", X"00", X"7c", 
  X"af", X"ab", X"00", X"80", X"24", X"42", X"00", X"01", 
  X"af", X"a2", X"00", X"7c", X"28", X"42", X"00", X"08", 
  X"14", X"40", X"00", X"07", X"25", X"29", X"00", X"08", 
  X"02", X"40", X"20", X"21", X"02", X"20", X"28", X"21", 
  X"0f", X"f0", X"06", X"a5", X"27", X"a6", X"00", X"78", 
  X"14", X"40", X"00", X"4b", X"27", X"a9", X"00", X"10", 
  X"32", X"8a", X"00", X"04", X"15", X"40", X"00", X"0c", 
  X"8f", X"a3", X"00", X"88", X"8f", X"a5", X"00", X"88", 
  X"02", X"a5", X"10", X"2a", X"00", X"a2", X"a8", X"0b", 
  X"8f", X"a2", X"00", X"8c", X"00", X"55", X"10", X"21", 
  X"af", X"a2", X"00", X"8c", X"8f", X"a2", X"00", X"80", 
  X"50", X"40", X"00", X"36", X"af", X"a0", X"00", X"7c", 
  X"0b", X"f0", X"0a", X"11", X"02", X"40", X"20", X"21", 
  X"00", X"75", X"80", X"23", X"1a", X"00", X"ff", X"f3", 
  X"24", X"16", X"00", X"10", X"2a", X"04", X"00", X"11", 
  X"8f", X"a3", X"00", X"80", X"14", X"80", X"00", X"15", 
  X"8f", X"a2", X"00", X"7c", X"24", X"42", X"00", X"01", 
  X"3c", X"04", X"bf", X"c0", X"24", X"84", X"5c", X"50", 
  X"24", X"63", X"00", X"10", X"af", X"a2", X"00", X"7c", 
  X"28", X"42", X"00", X"08", X"ad", X"24", X"00", X"00", 
  X"ad", X"36", X"00", X"04", X"10", X"40", X"00", X"03", 
  X"af", X"a3", X"00", X"80", X"0b", X"f0", X"09", X"fd", 
  X"25", X"29", X"00", X"08", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"14", X"40", X"00", X"24", 
  X"27", X"a9", X"00", X"10", X"0b", X"f0", X"09", X"e7", 
  X"26", X"10", X"ff", X"f0", X"24", X"42", X"00", X"01", 
  X"3c", X"05", X"bf", X"c0", X"24", X"a5", X"5c", X"50", 
  X"ad", X"30", X"00", X"04", X"af", X"a2", X"00", X"7c", 
  X"00", X"70", X"80", X"21", X"28", X"42", X"00", X"08", 
  X"ad", X"25", X"00", X"00", X"14", X"40", X"ff", X"d1", 
  X"af", X"b0", X"00", X"80", X"02", X"40", X"20", X"21", 
  X"02", X"20", X"28", X"21", X"0f", X"f0", X"06", X"a5", 
  X"27", X"a6", X"00", X"78", X"10", X"40", X"ff", X"cc", 
  X"8f", X"a5", X"00", X"88", X"0b", X"f0", X"0a", X"21", 
  X"96", X"22", X"00", X"0c", X"02", X"20", X"28", X"21", 
  X"0f", X"f0", X"06", X"a5", X"27", X"a6", X"00", X"78", 
  X"54", X"40", X"00", X"0c", X"96", X"22", X"00", X"0c", 
  X"af", X"a0", X"00", X"7c", X"0b", X"f0", X"07", X"25", 
  X"27", X"a9", X"00", X"10", X"8f", X"a2", X"00", X"80", 
  X"50", X"40", X"00", X"06", X"96", X"22", X"00", X"0c", 
  X"02", X"40", X"20", X"21", X"02", X"20", X"28", X"21", 
  X"0f", X"f0", X"06", X"a5", X"27", X"a6", X"00", X"78", 
  X"96", X"22", X"00", X"0c", X"30", X"42", X"00", X"40", 
  X"14", X"40", X"00", X"02", X"24", X"02", X"ff", X"ff", 
  X"8f", X"a2", X"00", X"8c", X"8f", X"bf", X"00", X"c4", 
  X"8f", X"be", X"00", X"c0", X"8f", X"b7", X"00", X"bc", 
  X"8f", X"b6", X"00", X"b8", X"8f", X"b5", X"00", X"b4", 
  X"8f", X"b4", X"00", X"b0", X"8f", X"b3", X"00", X"ac", 
  X"8f", X"b2", X"00", X"a8", X"8f", X"b1", X"00", X"a4", 
  X"8f", X"b0", X"00", X"a0", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"c8", X"00", X"80", X"18", X"21", 
  X"3c", X"04", X"00", X"00", X"8c", X"84", X"08", X"9c", 
  X"00", X"a0", X"10", X"21", X"00", X"c0", X"38", X"21", 
  X"00", X"60", X"28", X"21", X"0b", X"f0", X"06", X"e3", 
  X"00", X"40", X"30", X"21", X"94", X"a2", X"00", X"0c", 
  X"27", X"bd", X"fb", X"78", X"af", X"b0", X"04", X"78", 
  X"30", X"42", X"ff", X"fd", X"a7", X"a2", X"04", X"1c", 
  X"8c", X"a2", X"00", X"60", X"00", X"a0", X"80", X"21", 
  X"af", X"b2", X"04", X"80", X"af", X"a2", X"04", X"70", 
  X"94", X"a2", X"00", X"0e", X"af", X"b1", X"04", X"7c", 
  X"af", X"bf", X"04", X"84", X"a7", X"a2", X"04", X"1e", 
  X"8c", X"a2", X"00", X"1c", X"00", X"80", X"90", X"21", 
  X"af", X"a0", X"04", X"28", X"af", X"a2", X"04", X"2c", 
  X"8c", X"a2", X"00", X"24", X"27", X"a5", X"04", X"10", 
  X"af", X"a2", X"04", X"34", X"27", X"a2", X"00", X"10", 
  X"af", X"a2", X"04", X"10", X"af", X"a2", X"04", X"20", 
  X"24", X"02", X"04", X"00", X"af", X"a2", X"04", X"18", 
  X"0f", X"f0", X"06", X"e3", X"af", X"a2", X"04", X"24", 
  X"04", X"40", X"00", X"06", X"00", X"40", X"88", X"21", 
  X"02", X"40", X"20", X"21", X"0f", X"f0", X"0b", X"46", 
  X"27", X"a5", X"04", X"10", X"24", X"03", X"ff", X"ff", 
  X"00", X"62", X"88", X"0b", X"97", X"a2", X"04", X"1c", 
  X"30", X"42", X"00", X"40", X"10", X"40", X"00", X"05", 
  X"8f", X"bf", X"04", X"84", X"96", X"02", X"00", X"0c", 
  X"34", X"42", X"00", X"40", X"a6", X"02", X"00", X"0c", 
  X"8f", X"bf", X"04", X"84", X"02", X"20", X"10", X"21", 
  X"8f", X"b2", X"04", X"80", X"8f", X"b1", X"04", X"7c", 
  X"8f", X"b0", X"04", X"78", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"04", X"88", X"27", X"bd", X"ff", X"e0", 
  X"3c", X"02", X"00", X"00", X"af", X"b1", X"00", X"18", 
  X"00", X"80", X"88", X"21", X"8c", X"44", X"08", X"9c", 
  X"af", X"b0", X"00", X"14", X"af", X"bf", X"00", X"1c", 
  X"10", X"80", X"00", X"06", X"00", X"a0", X"80", X"21", 
  X"8c", X"82", X"00", X"38", X"54", X"40", X"00", X"04", 
  X"86", X"03", X"00", X"0c", X"0f", X"f0", X"0b", X"91", 
  X"00", X"00", X"00", X"00", X"86", X"03", X"00", X"0c", 
  X"30", X"62", X"ff", X"ff", X"30", X"44", X"00", X"08", 
  X"54", X"80", X"00", X"1b", X"8e", X"02", X"00", X"10", 
  X"30", X"44", X"00", X"10", X"14", X"80", X"00", X"04", 
  X"30", X"42", X"00", X"04", X"24", X"02", X"00", X"09", 
  X"0b", X"f0", X"0a", X"b3", X"ae", X"22", X"00", X"00", 
  X"50", X"40", X"00", X"10", X"96", X"02", X"00", X"0c", 
  X"8e", X"05", X"00", X"30", X"10", X"a0", X"00", X"06", 
  X"26", X"02", X"00", X"40", X"50", X"a2", X"00", X"04", 
  X"ae", X"00", X"00", X"30", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"20", X"20", X"21", X"ae", X"00", X"00", X"30", 
  X"96", X"02", X"00", X"0c", X"ae", X"00", X"00", X"04", 
  X"30", X"42", X"ff", X"db", X"a6", X"02", X"00", X"0c", 
  X"8e", X"02", X"00", X"10", X"ae", X"02", X"00", X"00", 
  X"96", X"02", X"00", X"0c", X"34", X"42", X"00", X"08", 
  X"a6", X"02", X"00", X"0c", X"8e", X"02", X"00", X"10", 
  X"54", X"40", X"00", X"09", X"96", X"02", X"00", X"0c", 
  X"96", X"03", X"00", X"0c", X"24", X"02", X"02", X"00", 
  X"30", X"63", X"02", X"80", X"10", X"62", X"00", X"03", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"0f", X"3e", 
  X"02", X"00", X"28", X"21", X"96", X"02", X"00", X"0c", 
  X"30", X"43", X"00", X"01", X"10", X"60", X"00", X"06", 
  X"30", X"43", X"00", X"02", X"8e", X"02", X"00", X"14", 
  X"ae", X"00", X"00", X"08", X"00", X"02", X"10", X"23", 
  X"0b", X"f0", X"0a", X"ac", X"ae", X"02", X"00", X"18", 
  X"14", X"60", X"00", X"02", X"00", X"00", X"10", X"21", 
  X"8e", X"02", X"00", X"14", X"ae", X"02", X"00", X"08", 
  X"8e", X"03", X"00", X"10", X"14", X"60", X"00", X"08", 
  X"00", X"00", X"10", X"21", X"86", X"03", X"00", X"0c", 
  X"30", X"64", X"00", X"80", X"10", X"80", X"00", X"05", 
  X"8f", X"bf", X"00", X"1c", X"34", X"63", X"00", X"40", 
  X"a6", X"03", X"00", X"0c", X"24", X"02", X"ff", X"ff", 
  X"8f", X"bf", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"84", X"a2", X"00", X"0c", 
  X"27", X"bd", X"ff", X"d8", X"af", X"b1", X"00", X"18", 
  X"30", X"43", X"00", X"08", X"af", X"b0", X"00", X"14", 
  X"af", X"bf", X"00", X"24", X"af", X"b3", X"00", X"20", 
  X"af", X"b2", X"00", X"1c", X"00", X"80", X"88", X"21", 
  X"14", X"60", X"00", X"5d", X"00", X"a0", X"80", X"21", 
  X"8c", X"a3", X"00", X"04", X"34", X"42", X"08", X"00", 
  X"1c", X"60", X"00", X"04", X"a4", X"a2", X"00", X"0c", 
  X"8c", X"a3", X"00", X"3c", X"58", X"60", X"00", X"73", 
  X"00", X"00", X"10", X"21", X"8e", X"03", X"00", X"28", 
  X"50", X"60", X"00", X"70", X"00", X"00", X"10", X"21", 
  X"30", X"42", X"10", X"00", X"8e", X"32", X"00", X"00", 
  X"10", X"40", X"00", X"03", X"ae", X"20", X"00", X"00", 
  X"0b", X"f0", X"0a", X"e9", X"8e", X"02", X"00", X"50", 
  X"8e", X"05", X"00", X"1c", X"02", X"20", X"20", X"21", 
  X"00", X"00", X"30", X"21", X"00", X"60", X"f8", X"09", 
  X"24", X"07", X"00", X"01", X"24", X"03", X"ff", X"ff", 
  X"54", X"43", X"00", X"0d", X"96", X"03", X"00", X"0c", 
  X"8e", X"23", X"00", X"00", X"50", X"60", X"00", X"0a", 
  X"96", X"03", X"00", X"0c", X"24", X"02", X"00", X"1d", 
  X"50", X"62", X"00", X"3b", X"ae", X"32", X"00", X"00", 
  X"24", X"02", X"00", X"16", X"54", X"62", X"00", X"49", 
  X"96", X"02", X"00", X"0c", X"0b", X"f0", X"0b", X"1e", 
  X"ae", X"32", X"00", X"00", X"96", X"03", X"00", X"0c", 
  X"30", X"63", X"00", X"04", X"50", X"60", X"00", X"09", 
  X"8e", X"03", X"00", X"28", X"8e", X"03", X"00", X"04", 
  X"00", X"43", X"10", X"23", X"8e", X"03", X"00", X"30", 
  X"50", X"60", X"00", X"04", X"8e", X"03", X"00", X"28", 
  X"8e", X"03", X"00", X"3c", X"00", X"43", X"10", X"23", 
  X"8e", X"03", X"00", X"28", X"8e", X"05", X"00", X"1c", 
  X"02", X"20", X"20", X"21", X"00", X"40", X"30", X"21", 
  X"00", X"60", X"f8", X"09", X"00", X"00", X"38", X"21", 
  X"24", X"03", X"ff", X"ff", X"14", X"43", X"00", X"09", 
  X"96", X"04", X"00", X"0c", X"8e", X"23", X"00", X"00", 
  X"50", X"60", X"00", X"07", X"24", X"03", X"f7", X"ff", 
  X"24", X"05", X"00", X"1d", X"10", X"65", X"00", X"03", 
  X"24", X"05", X"00", X"16", X"54", X"65", X"00", X"1c", 
  X"34", X"84", X"00", X"40", X"24", X"03", X"f7", X"ff", 
  X"00", X"83", X"20", X"24", X"8e", X"03", X"00", X"10", 
  X"7c", X"04", X"26", X"20", X"a6", X"04", X"00", X"0c", 
  X"30", X"84", X"10", X"00", X"ae", X"00", X"00", X"04", 
  X"10", X"80", X"00", X"08", X"ae", X"03", X"00", X"00", 
  X"24", X"03", X"ff", X"ff", X"54", X"43", X"00", X"05", 
  X"ae", X"02", X"00", X"50", X"8e", X"23", X"00", X"00", 
  X"54", X"60", X"00", X"03", X"8e", X"05", X"00", X"30", 
  X"ae", X"02", X"00", X"50", X"8e", X"05", X"00", X"30", 
  X"10", X"a0", X"00", X"07", X"ae", X"32", X"00", X"00", 
  X"26", X"02", X"00", X"40", X"50", X"a2", X"00", X"04", 
  X"ae", X"00", X"00", X"30", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"20", X"20", X"21", X"ae", X"00", X"00", X"30", 
  X"0b", X"f0", X"0b", X"3f", X"00", X"00", X"10", X"21", 
  X"0b", X"f0", X"0b", X"31", X"a6", X"04", X"00", X"0c", 
  X"8c", X"b2", X"00", X"10", X"52", X"40", X"00", X"1b", 
  X"00", X"00", X"10", X"21", X"8c", X"b3", X"00", X"00", 
  X"30", X"42", X"00", X"03", X"ac", X"b2", X"00", X"00", 
  X"02", X"72", X"98", X"23", X"14", X"40", X"00", X"02", 
  X"00", X"00", X"18", X"21", X"8c", X"a3", X"00", X"14", 
  X"0b", X"f0", X"0b", X"3b", X"ae", X"03", X"00", X"08", 
  X"96", X"02", X"00", X"0c", X"34", X"42", X"00", X"40", 
  X"a6", X"02", X"00", X"0c", X"0b", X"f0", X"0b", X"3f", 
  X"24", X"02", X"ff", X"ff", X"8e", X"05", X"00", X"1c", 
  X"02", X"20", X"20", X"21", X"02", X"40", X"30", X"21", 
  X"00", X"40", X"f8", X"09", X"02", X"60", X"38", X"21", 
  X"18", X"40", X"ff", X"f5", X"02", X"42", X"90", X"21", 
  X"02", X"62", X"98", X"23", X"5e", X"60", X"ff", X"f7", 
  X"8e", X"02", X"00", X"24", X"0b", X"f0", X"0b", X"3f", 
  X"00", X"00", X"10", X"21", X"8f", X"bf", X"00", X"24", 
  X"8f", X"b3", X"00", X"20", X"8f", X"b2", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b0", X"00", X"18", 
  X"af", X"bf", X"00", X"1c", X"10", X"80", X"00", X"07", 
  X"00", X"80", X"80", X"21", X"8c", X"82", X"00", X"38", 
  X"54", X"40", X"00", X"05", X"84", X"a2", X"00", X"0c", 
  X"0f", X"f0", X"0b", X"91", X"af", X"a5", X"00", X"10", 
  X"8f", X"a5", X"00", X"10", X"84", X"a2", X"00", X"0c", 
  X"10", X"40", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"02", X"00", X"20", X"21", X"8f", X"b0", X"00", X"18", 
  X"0b", X"f0", X"0a", X"bb", X"27", X"bd", X"00", X"20", 
  X"8f", X"b0", X"00", X"18", X"00", X"00", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"14", X"80", X"00", X"0b", X"00", X"80", X"28", X"21", 
  X"3c", X"02", X"00", X"00", X"8c", X"44", X"08", X"98", 
  X"3c", X"05", X"bf", X"c0", X"27", X"bd", X"ff", X"e8", 
  X"af", X"bf", X"00", X"14", X"0f", X"f0", X"0e", X"dc", 
  X"24", X"a5", X"2d", X"18", X"8f", X"bf", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"18", 
  X"3c", X"02", X"00", X"00", X"0b", X"f0", X"0b", X"46", 
  X"8c", X"44", X"08", X"9c", X"3c", X"05", X"bf", X"c0", 
  X"27", X"bd", X"ff", X"e8", X"af", X"bf", X"00", X"14", 
  X"0f", X"f0", X"0e", X"b4", X"24", X"a5", X"59", X"1c", 
  X"8f", X"bf", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"18", X"27", X"bd", X"ff", X"e0", 
  X"24", X"02", X"00", X"64", X"af", X"b1", X"00", X"14", 
  X"24", X"b1", X"ff", X"ff", X"72", X"22", X"88", X"02", 
  X"af", X"b2", X"00", X"18", X"00", X"a0", X"90", X"21", 
  X"af", X"b0", X"00", X"10", X"af", X"bf", X"00", X"1c", 
  X"0f", X"f0", X"0f", X"94", X"26", X"25", X"00", X"70", 
  X"10", X"40", X"00", X"08", X"00", X"40", X"80", X"21", 
  X"24", X"44", X"00", X"0c", X"ac", X"40", X"00", X"00", 
  X"ac", X"52", X"00", X"04", X"ac", X"44", X"00", X"08", 
  X"00", X"00", X"28", X"21", X"0f", X"f0", X"12", X"53", 
  X"26", X"26", X"00", X"64", X"8f", X"bf", X"00", X"1c", 
  X"02", X"00", X"10", X"21", X"8f", X"b2", X"00", X"18", 
  X"8f", X"b1", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"3c", X"02", X"00", X"00", X"0b", X"f0", X"0b", X"6b", 
  X"8c", X"44", X"08", X"98", X"8c", X"82", X"00", X"38", 
  X"27", X"bd", X"ff", X"d0", X"af", X"b1", X"00", X"18", 
  X"af", X"bf", X"00", X"2c", X"af", X"b5", X"00", X"28", 
  X"af", X"b4", X"00", X"24", X"af", X"b3", X"00", X"20", 
  X"af", X"b2", X"00", X"1c", X"af", X"b0", X"00", X"14", 
  X"14", X"40", X"00", X"51", X"00", X"80", X"88", X"21", 
  X"3c", X"02", X"bf", X"c0", X"24", X"42", X"2d", X"ac", 
  X"8c", X"90", X"00", X"04", X"ac", X"82", X"00", X"3c", 
  X"24", X"02", X"00", X"03", X"ac", X"82", X"02", X"e4", 
  X"24", X"82", X"02", X"ec", X"ac", X"82", X"02", X"e8", 
  X"3c", X"15", X"bf", X"c0", X"24", X"02", X"00", X"04", 
  X"3c", X"14", X"bf", X"c0", X"3c", X"13", X"bf", X"c0", 
  X"3c", X"12", X"bf", X"c0", X"ac", X"80", X"02", X"e0", 
  X"26", X"b5", X"50", X"a4", X"26", X"04", X"00", X"58", 
  X"26", X"94", X"50", X"f8", X"26", X"73", X"51", X"78", 
  X"26", X"52", X"51", X"c8", X"ae", X"00", X"00", X"00", 
  X"ae", X"00", X"00", X"04", X"ae", X"00", X"00", X"08", 
  X"a6", X"02", X"00", X"0c", X"ae", X"00", X"00", X"60", 
  X"a6", X"00", X"00", X"0e", X"ae", X"00", X"00", X"10", 
  X"ae", X"00", X"00", X"14", X"ae", X"00", X"00", X"18", 
  X"00", X"00", X"28", X"21", X"0f", X"f0", X"12", X"53", 
  X"24", X"06", X"00", X"08", X"ae", X"10", X"00", X"1c", 
  X"ae", X"15", X"00", X"20", X"ae", X"14", X"00", X"24", 
  X"ae", X"13", X"00", X"28", X"ae", X"12", X"00", X"2c", 
  X"8e", X"30", X"00", X"08", X"24", X"02", X"00", X"09", 
  X"00", X"00", X"28", X"21", X"a6", X"02", X"00", X"0c", 
  X"24", X"02", X"00", X"01", X"26", X"04", X"00", X"58", 
  X"ae", X"00", X"00", X"00", X"ae", X"00", X"00", X"04", 
  X"ae", X"00", X"00", X"08", X"ae", X"00", X"00", X"60", 
  X"a6", X"02", X"00", X"0e", X"ae", X"00", X"00", X"10", 
  X"ae", X"00", X"00", X"14", X"ae", X"00", X"00", X"18", 
  X"0f", X"f0", X"12", X"53", X"24", X"06", X"00", X"08", 
  X"ae", X"10", X"00", X"1c", X"ae", X"15", X"00", X"20", 
  X"ae", X"14", X"00", X"24", X"ae", X"13", X"00", X"28", 
  X"ae", X"12", X"00", X"2c", X"8e", X"30", X"00", X"0c", 
  X"24", X"02", X"00", X"12", X"00", X"00", X"28", X"21", 
  X"a6", X"02", X"00", X"0c", X"24", X"02", X"00", X"02", 
  X"ae", X"00", X"00", X"00", X"ae", X"00", X"00", X"04", 
  X"ae", X"00", X"00", X"08", X"ae", X"00", X"00", X"60", 
  X"a6", X"02", X"00", X"0e", X"ae", X"00", X"00", X"10", 
  X"ae", X"00", X"00", X"14", X"ae", X"00", X"00", X"18", 
  X"26", X"04", X"00", X"58", X"0f", X"f0", X"12", X"53", 
  X"24", X"06", X"00", X"08", X"24", X"02", X"00", X"01", 
  X"ae", X"10", X"00", X"1c", X"ae", X"15", X"00", X"20", 
  X"ae", X"14", X"00", X"24", X"ae", X"13", X"00", X"28", 
  X"ae", X"12", X"00", X"2c", X"ae", X"22", X"00", X"38", 
  X"8f", X"bf", X"00", X"2c", X"8f", X"b5", X"00", X"28", 
  X"8f", X"b4", X"00", X"24", X"8f", X"b3", X"00", X"20", 
  X"8f", X"b2", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"27", X"bd", X"ff", X"e0", 
  X"3c", X"02", X"00", X"00", X"af", X"b1", X"00", X"14", 
  X"8c", X"51", X"08", X"98", X"af", X"b2", X"00", X"18", 
  X"af", X"bf", X"00", X"1c", X"8e", X"22", X"00", X"38", 
  X"af", X"b0", X"00", X"10", X"14", X"40", X"00", X"03", 
  X"00", X"80", X"90", X"21", X"0f", X"f0", X"0b", X"91", 
  X"02", X"20", X"20", X"21", X"26", X"31", X"02", X"e0", 
  X"8e", X"30", X"00", X"08", X"8e", X"22", X"00", X"04", 
  X"24", X"42", X"ff", X"ff", X"04", X"42", X"00", X"06", 
  X"8e", X"22", X"00", X"00", X"86", X"03", X"00", X"0c", 
  X"50", X"60", X"00", X"10", X"24", X"02", X"ff", X"ff", 
  X"0b", X"f0", X"0c", X"04", X"26", X"10", X"00", X"64", 
  X"54", X"40", X"ff", X"f5", X"8e", X"31", X"00", X"00", 
  X"02", X"40", X"20", X"21", X"0f", X"f0", X"0b", X"73", 
  X"24", X"05", X"00", X"04", X"10", X"40", X"00", X"03", 
  X"ae", X"22", X"00", X"00", X"0b", X"f0", X"0c", X"02", 
  X"8e", X"31", X"00", X"00", X"24", X"02", X"00", X"0c", 
  X"ae", X"42", X"00", X"00", X"0b", X"f0", X"0c", X"2c", 
  X"00", X"00", X"10", X"21", X"a6", X"02", X"00", X"0e", 
  X"24", X"02", X"00", X"01", X"a6", X"02", X"00", X"0c", 
  X"ae", X"00", X"00", X"60", X"ae", X"00", X"00", X"00", 
  X"ae", X"00", X"00", X"08", X"ae", X"00", X"00", X"04", 
  X"ae", X"00", X"00", X"10", X"ae", X"00", X"00", X"14", 
  X"ae", X"00", X"00", X"18", X"26", X"04", X"00", X"58", 
  X"00", X"00", X"28", X"21", X"0f", X"f0", X"12", X"53", 
  X"24", X"06", X"00", X"08", X"ae", X"00", X"00", X"30", 
  X"ae", X"00", X"00", X"34", X"ae", X"00", X"00", X"44", 
  X"ae", X"00", X"00", X"48", X"02", X"00", X"10", X"21", 
  X"8f", X"bf", X"00", X"1c", X"8f", X"b2", X"00", X"18", 
  X"8f", X"b1", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"84", X"c2", X"00", X"0c", X"27", X"bd", X"ff", X"c8", 
  X"af", X"b3", X"00", X"28", X"30", X"43", X"20", X"00", 
  X"af", X"b2", X"00", X"24", X"af", X"b0", X"00", X"1c", 
  X"af", X"bf", X"00", X"34", X"af", X"b5", X"00", X"30", 
  X"af", X"b4", X"00", X"2c", X"af", X"b1", X"00", X"20", 
  X"00", X"80", X"98", X"21", X"00", X"a0", X"90", X"21", 
  X"14", X"60", X"00", X"06", X"00", X"c0", X"80", X"21", 
  X"34", X"42", X"20", X"00", X"a4", X"c2", X"00", X"0c", 
  X"8c", X"c2", X"00", X"60", X"34", X"42", X"20", X"00", 
  X"ac", X"c2", X"00", X"60", X"0f", X"f0", X"0f", X"2a", 
  X"00", X"00", X"00", X"00", X"24", X"03", X"00", X"01", 
  X"14", X"43", X"00", X"07", X"02", X"60", X"20", X"21", 
  X"26", X"42", X"ff", X"ff", X"2c", X"42", X"00", X"ff", 
  X"10", X"40", X"00", X"03", X"24", X"02", X"00", X"01", 
  X"0b", X"f0", X"0c", X"5b", X"a3", X"b2", X"00", X"10", 
  X"27", X"a5", X"00", X"10", X"02", X"40", X"30", X"21", 
  X"0f", X"f0", X"15", X"8f", X"26", X"07", X"00", X"58", 
  X"24", X"03", X"ff", X"ff", X"14", X"43", X"00", X"06", 
  X"27", X"b1", X"00", X"10", X"96", X"02", X"00", X"0c", 
  X"34", X"42", X"00", X"40", X"0b", X"f0", X"0c", X"85", 
  X"a6", X"02", X"00", X"0c", X"27", X"b1", X"00", X"10", 
  X"02", X"22", X"a0", X"21", X"24", X"15", X"00", X"0a", 
  X"12", X"34", X"00", X"27", X"02", X"40", X"10", X"21", 
  X"8e", X"03", X"00", X"08", X"24", X"63", X"ff", X"ff", 
  X"04", X"61", X"00", X"1a", X"ae", X"03", X"00", X"08", 
  X"8e", X"02", X"00", X"18", X"00", X"62", X"18", X"2a", 
  X"54", X"60", X"00", X"0d", X"92", X"25", X"00", X"00", 
  X"8e", X"02", X"00", X"00", X"92", X"23", X"00", X"00", 
  X"a0", X"43", X"00", X"00", X"8e", X"03", X"00", X"00", 
  X"90", X"62", X"00", X"00", X"10", X"55", X"00", X"03", 
  X"24", X"63", X"00", X"01", X"0b", X"f0", X"0c", X"83", 
  X"ae", X"03", X"00", X"00", X"02", X"60", X"20", X"21", 
  X"0b", X"f0", X"0c", X"75", X"24", X"05", X"00", X"0a", 
  X"02", X"60", X"20", X"21", X"0f", X"f0", X"15", X"37", 
  X"02", X"00", X"30", X"21", X"24", X"42", X"00", X"01", 
  X"2c", X"43", X"00", X"01", X"10", X"60", X"ff", X"e4", 
  X"26", X"31", X"00", X"01", X"0b", X"f0", X"0c", X"86", 
  X"24", X"02", X"ff", X"ff", X"8e", X"02", X"00", X"00", 
  X"92", X"23", X"00", X"00", X"a0", X"43", X"00", X"00", 
  X"8e", X"02", X"00", X"00", X"24", X"42", X"00", X"01", 
  X"ae", X"02", X"00", X"00", X"0b", X"f0", X"0c", X"5e", 
  X"26", X"31", X"00", X"01", X"24", X"02", X"ff", X"ff", 
  X"8f", X"bf", X"00", X"34", X"8f", X"b5", X"00", X"30", 
  X"8f", X"b4", X"00", X"2c", X"8f", X"b3", X"00", X"28", 
  X"8f", X"b2", X"00", X"24", X"8f", X"b1", X"00", X"20", 
  X"8f", X"b0", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"27", X"bd", X"ff", X"e0", 
  X"3c", X"02", X"00", X"00", X"af", X"b0", X"00", X"10", 
  X"8c", X"50", X"08", X"9c", X"af", X"b2", X"00", X"18", 
  X"af", X"b1", X"00", X"14", X"af", X"bf", X"00", X"1c", 
  X"00", X"80", X"90", X"21", X"12", X"00", X"00", X"06", 
  X"00", X"a0", X"88", X"21", X"8e", X"02", X"00", X"38", 
  X"14", X"40", X"00", X"04", X"8f", X"bf", X"00", X"1c", 
  X"0f", X"f0", X"0b", X"91", X"02", X"00", X"20", X"21", 
  X"8f", X"bf", X"00", X"1c", X"02", X"00", X"20", X"21", 
  X"02", X"40", X"28", X"21", X"8f", X"b0", X"00", X"10", 
  X"8f", X"b2", X"00", X"18", X"02", X"20", X"30", X"21", 
  X"8f", X"b1", X"00", X"14", X"0b", X"f0", X"0c", X"32", 
  X"27", X"bd", X"00", X"20", X"27", X"bd", X"ff", X"d8", 
  X"af", X"b2", X"00", X"1c", X"3c", X"12", X"00", X"00", 
  X"26", X"52", X"04", X"90", X"af", X"b3", X"00", X"20", 
  X"af", X"b1", X"00", X"18", X"af", X"b0", X"00", X"14", 
  X"00", X"a0", X"88", X"21", X"af", X"bf", X"00", X"24", 
  X"0f", X"f0", X"12", X"9e", X"00", X"80", X"80", X"21", 
  X"8e", X"42", X"00", X"08", X"24", X"13", X"ff", X"fc", 
  X"8c", X"42", X"00", X"04", X"02", X"62", X"98", X"24", 
  X"02", X"71", X"88", X"23", X"26", X"31", X"0f", X"ef", 
  X"00", X"11", X"8b", X"02", X"26", X"31", X"ff", X"ff", 
  X"00", X"11", X"8b", X"00", X"2a", X"22", X"10", X"00", 
  X"10", X"40", X"00", X"05", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"12", X"a0", X"02", X"00", X"20", X"21", 
  X"0b", X"f0", X"0c", X"e6", X"00", X"00", X"10", X"21", 
  X"0f", X"f0", X"14", X"15", X"00", X"00", X"28", X"21", 
  X"8e", X"43", X"00", X"08", X"00", X"73", X"18", X"21", 
  X"14", X"43", X"ff", X"f7", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"14", X"15", X"00", X"11", X"28", X"23", 
  X"24", X"03", X"ff", X"ff", X"54", X"43", X"00", X"10", 
  X"8e", X"42", X"00", X"08", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"14", X"15", X"00", X"00", X"28", X"21", 
  X"8e", X"43", X"00", X"08", X"00", X"43", X"20", X"23", 
  X"28", X"85", X"00", X"10", X"14", X"a0", X"ff", X"ea", 
  X"3c", X"05", X"00", X"00", X"8c", X"a5", X"08", X"a4", 
  X"34", X"84", X"00", X"01", X"ac", X"64", X"00", X"04", 
  X"00", X"45", X"10", X"23", X"3c", X"05", X"00", X"00", 
  X"0b", X"f0", X"0c", X"be", X"ac", X"a2", X"08", X"cc", 
  X"02", X"71", X"98", X"23", X"36", X"73", X"00", X"01", 
  X"ac", X"53", X"00", X"04", X"3c", X"02", X"00", X"00", 
  X"8c", X"43", X"08", X"cc", X"02", X"00", X"20", X"21", 
  X"00", X"71", X"88", X"23", X"0f", X"f0", X"12", X"a0", 
  X"ac", X"51", X"08", X"cc", X"24", X"02", X"00", X"01", 
  X"8f", X"bf", X"00", X"24", X"8f", X"b3", X"00", X"20", 
  X"8f", X"b2", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"27", X"bd", X"ff", X"e0", 
  X"af", X"b1", X"00", X"18", X"af", X"bf", X"00", X"1c", 
  X"af", X"b0", X"00", X"14", X"10", X"a0", X"00", X"96", 
  X"00", X"a0", X"88", X"21", X"0f", X"f0", X"12", X"9e", 
  X"00", X"80", X"80", X"21", X"8e", X"28", X"ff", X"fc", 
  X"24", X"03", X"ff", X"fe", X"26", X"22", X"ff", X"f8", 
  X"01", X"03", X"18", X"24", X"00", X"43", X"38", X"21", 
  X"8c", X"e4", X"00", X"04", X"3c", X"06", X"00", X"00", 
  X"24", X"05", X"ff", X"fc", X"24", X"c6", X"04", X"90", 
  X"00", X"a4", X"20", X"24", X"8c", X"c5", X"00", X"08", 
  X"14", X"e5", X"00", X"19", X"31", X"08", X"00", X"01", 
  X"15", X"00", X"00", X"08", X"00", X"83", X"18", X"21", 
  X"8e", X"24", X"ff", X"f8", X"00", X"44", X"10", X"23", 
  X"8c", X"45", X"00", X"08", X"00", X"64", X"18", X"21", 
  X"8c", X"44", X"00", X"0c", X"ac", X"a4", X"00", X"0c", 
  X"ac", X"85", X"00", X"08", X"34", X"64", X"00", X"01", 
  X"ac", X"44", X"00", X"04", X"ac", X"c2", X"00", X"08", 
  X"3c", X"02", X"00", X"00", X"8c", X"44", X"08", X"a8", 
  X"00", X"64", X"18", X"2b", X"14", X"60", X"00", X"04", 
  X"3c", X"02", X"00", X"00", X"8c", X"45", X"0d", X"5c", 
  X"0f", X"f0", X"0c", X"a7", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"12", X"a0", X"02", X"00", X"20", X"21", 
  X"0b", X"f0", X"0d", X"89", X"8f", X"bf", X"00", X"1c", 
  X"ac", X"e4", X"00", X"04", X"15", X"00", X"00", X"0c", 
  X"00", X"00", X"28", X"21", X"8e", X"28", X"ff", X"f8", 
  X"3c", X"09", X"00", X"00", X"25", X"29", X"04", X"98", 
  X"00", X"48", X"10", X"23", X"00", X"68", X"18", X"21", 
  X"8c", X"48", X"00", X"08", X"51", X"09", X"00", X"04", 
  X"24", X"05", X"00", X"01", X"8c", X"49", X"00", X"0c", 
  X"ad", X"09", X"00", X"0c", X"ad", X"28", X"00", X"08", 
  X"00", X"e4", X"40", X"21", X"8d", X"08", X"00", X"04", 
  X"31", X"08", X"00", X"01", X"55", X"00", X"00", X"12", 
  X"34", X"64", X"00", X"01", X"00", X"64", X"18", X"21", 
  X"14", X"a0", X"00", X"0b", X"8c", X"e4", X"00", X"08", 
  X"3c", X"08", X"00", X"00", X"25", X"08", X"04", X"98", 
  X"54", X"88", X"00", X"08", X"8c", X"e7", X"00", X"0c", 
  X"ac", X"c2", X"00", X"14", X"ac", X"c2", X"00", X"10", 
  X"24", X"05", X"00", X"01", X"ac", X"44", X"00", X"0c", 
  X"0b", X"f0", X"0d", X"3d", X"ac", X"44", X"00", X"08", 
  X"8c", X"e7", X"00", X"0c", X"ac", X"87", X"00", X"0c", 
  X"ac", X"e4", X"00", X"08", X"34", X"64", X"00", X"01", 
  X"ac", X"44", X"00", X"04", X"00", X"43", X"20", X"21", 
  X"14", X"a0", X"ff", X"d5", X"ac", X"83", X"00", X"00", 
  X"2c", X"64", X"02", X"00", X"10", X"80", X"00", X"10", 
  X"00", X"03", X"2a", X"42", X"00", X"03", X"18", X"c2", 
  X"00", X"03", X"20", X"83", X"24", X"05", X"00", X"01", 
  X"00", X"85", X"20", X"04", X"8c", X"c5", X"00", X"04", 
  X"00", X"03", X"18", X"c0", X"00", X"85", X"20", X"25", 
  X"ac", X"c4", X"00", X"04", X"00", X"c3", X"30", X"21", 
  X"8c", X"c3", X"00", X"08", X"ac", X"46", X"00", X"0c", 
  X"ac", X"43", X"00", X"08", X"ac", X"c2", X"00", X"08", 
  X"0b", X"f0", X"0d", X"16", X"ac", X"62", X"00", X"0c", 
  X"2c", X"a4", X"00", X"05", X"10", X"80", X"00", X"04", 
  X"2c", X"a4", X"00", X"15", X"00", X"03", X"29", X"82", 
  X"0b", X"f0", X"0d", X"6c", X"24", X"a5", X"00", X"38", 
  X"10", X"80", X"00", X"03", X"2c", X"a4", X"00", X"55", 
  X"0b", X"f0", X"0d", X"6c", X"24", X"a5", X"00", X"5b", 
  X"10", X"80", X"00", X"04", X"2c", X"a4", X"01", X"55", 
  X"00", X"03", X"2b", X"02", X"0b", X"f0", X"0d", X"6c", 
  X"24", X"a5", X"00", X"6e", X"10", X"80", X"00", X"04", 
  X"2c", X"a4", X"05", X"55", X"00", X"03", X"2b", X"c2", 
  X"0b", X"f0", X"0d", X"6c", X"24", X"a5", X"00", X"77", 
  X"10", X"80", X"00", X"03", X"24", X"05", X"00", X"7e", 
  X"00", X"03", X"2c", X"82", X"24", X"a5", X"00", X"7c", 
  X"00", X"05", X"20", X"c0", X"00", X"c4", X"20", X"21", 
  X"8c", X"87", X"00", X"08", X"50", X"e4", X"00", X"04", 
  X"24", X"03", X"00", X"01", X"00", X"e0", X"28", X"21", 
  X"0b", X"f0", X"0d", X"7d", X"24", X"07", X"ff", X"fc", 
  X"00", X"05", X"28", X"83", X"00", X"a3", X"28", X"04", 
  X"8c", X"c3", X"00", X"04", X"00", X"a3", X"28", X"25", 
  X"ac", X"c5", X"00", X"04", X"0b", X"f0", X"0d", X"83", 
  X"00", X"e0", X"28", X"21", X"50", X"a4", X"00", X"07", 
  X"8c", X"a7", X"00", X"0c", X"8c", X"a6", X"00", X"04", 
  X"00", X"e6", X"30", X"24", X"00", X"66", X"30", X"2b", 
  X"54", X"c0", X"ff", X"fa", X"8c", X"a5", X"00", X"08", 
  X"8c", X"a7", X"00", X"0c", X"ac", X"47", X"00", X"0c", 
  X"ac", X"45", X"00", X"08", X"ac", X"e2", X"00", X"08", 
  X"0b", X"f0", X"0d", X"16", X"ac", X"a2", X"00", X"0c", 
  X"8f", X"bf", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"8c", X"c2", X"00", X"08", 
  X"27", X"bd", X"ff", X"c0", X"af", X"b4", X"00", X"28", 
  X"af", X"bf", X"00", X"3c", X"af", X"be", X"00", X"38", 
  X"af", X"b7", X"00", X"34", X"af", X"b6", X"00", X"30", 
  X"af", X"b5", X"00", X"2c", X"af", X"b3", X"00", X"24", 
  X"af", X"b2", X"00", X"20", X"af", X"b1", X"00", X"1c", 
  X"af", X"b0", X"00", X"18", X"14", X"40", X"00", X"03", 
  X"00", X"c0", X"a0", X"21", X"0b", X"f0", X"0e", X"a8", 
  X"00", X"00", X"10", X"21", X"94", X"a2", X"00", X"0c", 
  X"00", X"80", X"98", X"21", X"30", X"42", X"00", X"08", 
  X"10", X"40", X"00", X"0c", X"00", X"a0", X"80", X"21", 
  X"8c", X"a2", X"00", X"10", X"10", X"40", X"00", X"0a", 
  X"02", X"60", X"20", X"21", X"96", X"02", X"00", X"0c", 
  X"30", X"43", X"00", X"02", X"10", X"60", X"00", X"21", 
  X"8e", X"92", X"00", X"00", X"00", X"00", X"a8", X"21", 
  X"00", X"00", X"88", X"21", X"0b", X"f0", X"0d", X"c3", 
  X"24", X"16", X"04", X"00", X"02", X"60", X"20", X"21", 
  X"0f", X"f0", X"0a", X"69", X"02", X"00", X"28", X"21", 
  X"50", X"40", X"ff", X"f5", X"96", X"02", X"00", X"0c", 
  X"0b", X"f0", X"0e", X"a8", X"24", X"02", X"ff", X"ff", 
  X"02", X"c0", X"18", X"21", X"8e", X"02", X"00", X"24", 
  X"8e", X"05", X"00", X"1c", X"02", X"27", X"18", X"0b", 
  X"02", X"60", X"20", X"21", X"02", X"a0", X"30", X"21", 
  X"00", X"40", X"f8", X"09", X"00", X"60", X"38", X"21", 
  X"18", X"40", X"00", X"e7", X"02", X"a2", X"a8", X"21", 
  X"8e", X"83", X"00", X"08", X"02", X"22", X"88", X"23", 
  X"00", X"62", X"10", X"23", X"10", X"40", X"ff", X"d9", 
  X"ae", X"82", X"00", X"08", X"56", X"20", X"ff", X"f0", 
  X"2e", X"27", X"04", X"01", X"8e", X"55", X"00", X"00", 
  X"8e", X"51", X"00", X"04", X"0b", X"f0", X"0d", X"c3", 
  X"26", X"52", X"00", X"08", X"30", X"42", X"00", X"01", 
  X"10", X"40", X"00", X"05", X"00", X"00", X"a8", X"21", 
  X"00", X"00", X"b8", X"21", X"00", X"00", X"18", X"21", 
  X"0b", X"f0", X"0e", X"76", X"00", X"00", X"b0", X"21", 
  X"00", X"00", X"b8", X"21", X"56", X"e0", X"00", X"05", 
  X"96", X"02", X"00", X"0c", X"8e", X"55", X"00", X"00", 
  X"8e", X"57", X"00", X"04", X"0b", X"f0", X"0d", X"d1", 
  X"26", X"52", X"00", X"08", X"8e", X"11", X"00", X"08", 
  X"30", X"45", X"02", X"00", X"10", X"a0", X"00", X"46", 
  X"8e", X"04", X"00", X"00", X"02", X"f1", X"28", X"2b", 
  X"54", X"a0", X"00", X"37", X"02", X"f1", X"10", X"2b", 
  X"30", X"45", X"04", X"80", X"50", X"a0", X"00", X"34", 
  X"02", X"f1", X"10", X"2b", X"8e", X"07", X"00", X"14", 
  X"24", X"03", X"00", X"03", X"8e", X"05", X"00", X"10", 
  X"70", X"67", X"38", X"02", X"30", X"42", X"04", X"00", 
  X"00", X"85", X"b0", X"23", X"00", X"07", X"27", X"c2", 
  X"00", X"87", X"38", X"21", X"26", X"c4", X"00", X"01", 
  X"00", X"97", X"20", X"21", X"00", X"07", X"f0", X"43", 
  X"03", X"c4", X"30", X"2b", X"00", X"86", X"f0", X"0b", 
  X"10", X"40", X"00", X"0f", X"02", X"60", X"20", X"21", 
  X"0f", X"f0", X"0f", X"94", X"03", X"c0", X"28", X"21", 
  X"10", X"40", X"00", X"15", X"00", X"40", X"88", X"21", 
  X"8e", X"05", X"00", X"10", X"00", X"40", X"20", X"21", 
  X"0f", X"f0", X"11", X"4e", X"02", X"c0", X"30", X"21", 
  X"96", X"02", X"00", X"0c", X"24", X"03", X"fb", X"7f", 
  X"00", X"43", X"10", X"24", X"34", X"42", X"00", X"80", 
  X"0b", X"f0", X"0e", X"0b", X"a6", X"02", X"00", X"0c", 
  X"0f", X"f0", X"12", X"a2", X"03", X"c0", X"30", X"21", 
  X"14", X"40", X"00", X"0a", X"00", X"40", X"88", X"21", 
  X"8e", X"05", X"00", X"10", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"60", X"20", X"21", X"96", X"02", X"00", X"0c", 
  X"30", X"42", X"ff", X"7f", X"a6", X"02", X"00", X"0c", 
  X"24", X"02", X"00", X"0c", X"0b", X"f0", X"0e", X"a4", 
  X"ae", X"62", X"00", X"00", X"ae", X"11", X"00", X"10", 
  X"02", X"36", X"88", X"21", X"03", X"d6", X"b0", X"23", 
  X"ae", X"11", X"00", X"00", X"ae", X"1e", X"00", X"14", 
  X"02", X"e0", X"88", X"21", X"ae", X"16", X"00", X"08", 
  X"02", X"f1", X"10", X"2b", X"8e", X"04", X"00", X"00", 
  X"02", X"e2", X"88", X"0b", X"02", X"20", X"30", X"21", 
  X"0f", X"f0", X"12", X"35", X"02", X"a0", X"28", X"21", 
  X"8e", X"02", X"00", X"08", X"00", X"51", X"10", X"23", 
  X"ae", X"02", X"00", X"08", X"8e", X"02", X"00", X"00", 
  X"00", X"51", X"88", X"21", X"ae", X"11", X"00", X"00", 
  X"0b", X"f0", X"0e", X"49", X"02", X"e0", X"88", X"21", 
  X"8e", X"02", X"00", X"10", X"00", X"44", X"10", X"2b", 
  X"50", X"40", X"00", X"11", X"8e", X"07", X"00", X"14", 
  X"02", X"37", X"10", X"2b", X"50", X"40", X"00", X"0e", 
  X"8e", X"07", X"00", X"14", X"02", X"a0", X"28", X"21", 
  X"0f", X"f0", X"12", X"35", X"02", X"20", X"30", X"21", 
  X"8e", X"02", X"00", X"00", X"02", X"60", X"20", X"21", 
  X"02", X"00", X"28", X"21", X"00", X"51", X"10", X"21", 
  X"0f", X"f0", X"0b", X"46", X"ae", X"02", X"00", X"00", 
  X"50", X"40", X"00", X"19", X"8e", X"82", X"00", X"08", 
  X"0b", X"f0", X"0e", X"a5", X"96", X"02", X"00", X"0c", 
  X"02", X"e7", X"10", X"2b", X"14", X"40", X"00", X"0a", 
  X"02", X"a0", X"28", X"21", X"8e", X"02", X"00", X"24", 
  X"8e", X"05", X"00", X"1c", X"02", X"60", X"20", X"21", 
  X"00", X"40", X"f8", X"09", X"02", X"a0", X"30", X"21", 
  X"1c", X"40", X"00", X"0c", X"00", X"40", X"88", X"21", 
  X"0b", X"f0", X"0e", X"a5", X"96", X"02", X"00", X"0c", 
  X"0f", X"f0", X"12", X"35", X"02", X"e0", X"30", X"21", 
  X"8e", X"02", X"00", X"08", X"02", X"e0", X"88", X"21", 
  X"00", X"57", X"10", X"23", X"ae", X"02", X"00", X"08", 
  X"8e", X"02", X"00", X"00", X"00", X"57", X"10", X"21", 
  X"ae", X"02", X"00", X"00", X"8e", X"82", X"00", X"08", 
  X"02", X"b1", X"a8", X"21", X"02", X"f1", X"b8", X"23", 
  X"00", X"51", X"88", X"23", X"16", X"20", X"ff", X"83", 
  X"ae", X"91", X"00", X"08", X"0b", X"f0", X"0e", X"a8", 
  X"00", X"00", X"10", X"21", X"10", X"60", X"00", X"2b", 
  X"02", X"c0", X"20", X"21", X"02", X"b7", X"f0", X"2b", 
  X"02", X"a0", X"10", X"21", X"02", X"fe", X"10", X"0a", 
  X"00", X"40", X"f0", X"21", X"8e", X"04", X"00", X"00", 
  X"8e", X"02", X"00", X"10", X"8e", X"11", X"00", X"08", 
  X"00", X"44", X"10", X"2b", X"10", X"40", X"00", X"2a", 
  X"8e", X"07", X"00", X"14", X"02", X"27", X"88", X"21", 
  X"02", X"3e", X"10", X"2a", X"10", X"40", X"00", X"27", 
  X"03", X"c7", X"10", X"2a", X"02", X"c0", X"28", X"21", 
  X"02", X"20", X"30", X"21", X"0f", X"f0", X"12", X"35", 
  X"af", X"a3", X"00", X"10", X"8e", X"02", X"00", X"00", 
  X"02", X"60", X"20", X"21", X"02", X"00", X"28", X"21", 
  X"00", X"51", X"10", X"21", X"0f", X"f0", X"0b", X"46", 
  X"ae", X"02", X"00", X"00", X"14", X"40", X"00", X"38", 
  X"8f", X"a3", X"00", X"10", X"02", X"f1", X"b8", X"23", 
  X"12", X"e0", X"00", X"31", X"02", X"60", X"20", X"21", 
  X"8e", X"82", X"00", X"08", X"02", X"d1", X"b0", X"21", 
  X"02", X"b1", X"a8", X"23", X"00", X"51", X"88", X"23", 
  X"12", X"20", X"ff", X"26", X"ae", X"91", X"00", X"08", 
  X"16", X"a0", X"ff", X"da", X"00", X"00", X"00", X"00", 
  X"8e", X"56", X"00", X"00", X"8e", X"55", X"00", X"04", 
  X"00", X"00", X"18", X"21", X"0b", X"f0", X"0e", X"76", 
  X"26", X"52", X"00", X"08", X"24", X"05", X"00", X"0a", 
  X"0f", X"f0", X"11", X"41", X"02", X"a0", X"30", X"21", 
  X"50", X"40", X"00", X"03", X"26", X"b7", X"00", X"01", 
  X"24", X"57", X"00", X"01", X"02", X"f6", X"b8", X"23", 
  X"0b", X"f0", X"0e", X"53", X"24", X"03", X"00", X"01", 
  X"03", X"c7", X"10", X"2a", X"14", X"40", X"00", X"0c", 
  X"02", X"c0", X"28", X"21", X"8e", X"02", X"00", X"24", 
  X"8e", X"05", X"00", X"1c", X"02", X"60", X"20", X"21", 
  X"af", X"a3", X"00", X"10", X"00", X"40", X"f8", X"09", 
  X"02", X"c0", X"30", X"21", X"00", X"40", X"88", X"21", 
  X"1c", X"40", X"ff", X"dc", X"8f", X"a3", X"00", X"10", 
  X"0b", X"f0", X"0e", X"a5", X"96", X"02", X"00", X"0c", 
  X"03", X"c0", X"30", X"21", X"0f", X"f0", X"12", X"35", 
  X"af", X"a3", X"00", X"10", X"8e", X"02", X"00", X"08", 
  X"03", X"c0", X"88", X"21", X"8f", X"a3", X"00", X"10", 
  X"00", X"5e", X"10", X"23", X"ae", X"02", X"00", X"08", 
  X"8e", X"02", X"00", X"00", X"00", X"5e", X"10", X"21", 
  X"0b", X"f0", X"0e", X"6d", X"ae", X"02", X"00", X"00", 
  X"0f", X"f0", X"0b", X"46", X"02", X"00", X"28", X"21", 
  X"10", X"40", X"ff", X"cd", X"00", X"00", X"18", X"21", 
  X"96", X"02", X"00", X"0c", X"34", X"42", X"00", X"40", 
  X"a6", X"02", X"00", X"0c", X"24", X"02", X"ff", X"ff", 
  X"8f", X"bf", X"00", X"3c", X"8f", X"be", X"00", X"38", 
  X"8f", X"b7", X"00", X"34", X"8f", X"b6", X"00", X"30", 
  X"8f", X"b5", X"00", X"2c", X"8f", X"b4", X"00", X"28", 
  X"8f", X"b3", X"00", X"24", X"8f", X"b2", X"00", X"20", 
  X"8f", X"b1", X"00", X"1c", X"8f", X"b0", X"00", X"18", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"40", 
  X"27", X"bd", X"ff", X"d0", X"af", X"b5", X"00", X"28", 
  X"af", X"b4", X"00", X"24", X"af", X"b2", X"00", X"1c", 
  X"af", X"b0", X"00", X"14", X"af", X"bf", X"00", X"2c", 
  X"af", X"b3", X"00", X"20", X"af", X"b1", X"00", X"18", 
  X"00", X"a0", X"a0", X"21", X"24", X"90", X"02", X"e0", 
  X"00", X"00", X"90", X"21", X"24", X"15", X"ff", X"ff", 
  X"12", X"00", X"00", X"12", X"8f", X"bf", X"00", X"2c", 
  X"8e", X"11", X"00", X"08", X"8e", X"13", X"00", X"04", 
  X"26", X"73", X"ff", X"ff", X"06", X"62", X"ff", X"fa", 
  X"8e", X"10", X"00", X"00", X"96", X"22", X"00", X"0c", 
  X"2c", X"42", X"00", X"02", X"54", X"40", X"ff", X"fa", 
  X"26", X"31", X"00", X"64", X"86", X"22", X"00", X"0e", 
  X"50", X"55", X"ff", X"f7", X"26", X"31", X"00", X"64", 
  X"02", X"80", X"f8", X"09", X"02", X"20", X"20", X"21", 
  X"02", X"42", X"90", X"25", X"0b", X"f0", X"0e", X"c4", 
  X"26", X"31", X"00", X"64", X"02", X"40", X"10", X"21", 
  X"8f", X"b5", X"00", X"28", X"8f", X"b4", X"00", X"24", 
  X"8f", X"b3", X"00", X"20", X"8f", X"b2", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"27", X"bd", X"ff", X"d0", X"af", X"b6", X"00", X"28", 
  X"af", X"b5", X"00", X"24", X"af", X"b4", X"00", X"20", 
  X"af", X"b2", X"00", X"18", X"af", X"b0", X"00", X"10", 
  X"af", X"bf", X"00", X"2c", X"af", X"b3", X"00", X"1c", 
  X"af", X"b1", X"00", X"14", X"00", X"80", X"a0", X"21", 
  X"00", X"a0", X"a8", X"21", X"24", X"90", X"02", X"e0", 
  X"00", X"00", X"90", X"21", X"24", X"16", X"ff", X"ff", 
  X"12", X"00", X"00", X"12", X"8f", X"bf", X"00", X"2c", 
  X"8e", X"11", X"00", X"08", X"8e", X"13", X"00", X"04", 
  X"26", X"73", X"ff", X"ff", X"06", X"62", X"ff", X"fa", 
  X"8e", X"10", X"00", X"00", X"96", X"22", X"00", X"0c", 
  X"2c", X"42", X"00", X"02", X"54", X"40", X"ff", X"fa", 
  X"26", X"31", X"00", X"64", X"86", X"22", X"00", X"0e", 
  X"10", X"56", X"00", X"04", X"02", X"80", X"20", X"21", 
  X"02", X"a0", X"f8", X"09", X"02", X"20", X"28", X"21", 
  X"02", X"42", X"90", X"25", X"0b", X"f0", X"0e", X"ee", 
  X"26", X"31", X"00", X"64", X"02", X"40", X"10", X"21", 
  X"8f", X"b6", X"00", X"28", X"8f", X"b5", X"00", X"24", 
  X"8f", X"b4", X"00", X"20", X"8f", X"b3", X"00", X"1c", 
  X"8f", X"b2", X"00", X"18", X"8f", X"b1", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"27", X"bd", X"ff", X"e0", 
  X"af", X"b1", X"00", X"18", X"af", X"b0", X"00", X"14", 
  X"af", X"bf", X"00", X"1c", X"00", X"c0", X"80", X"21", 
  X"14", X"c0", X"00", X"03", X"3c", X"11", X"bf", X"c0", 
  X"0b", X"f0", X"0f", X"22", X"26", X"22", X"5c", X"f8", 
  X"3c", X"05", X"bf", X"c0", X"00", X"c0", X"20", X"21", 
  X"0f", X"f0", X"14", X"7a", X"24", X"a5", X"5c", X"fc", 
  X"10", X"40", X"00", X"0d", X"26", X"22", X"5c", X"f8", 
  X"02", X"00", X"20", X"21", X"0f", X"f0", X"14", X"7a", 
  X"26", X"25", X"5c", X"f8", X"10", X"40", X"00", X"08", 
  X"26", X"22", X"5c", X"f8", X"3c", X"05", X"bf", X"c0", 
  X"02", X"00", X"20", X"21", X"0f", X"f0", X"14", X"7a", 
  X"24", X"a5", X"5c", X"ac", X"26", X"31", X"5c", X"f8", 
  X"00", X"02", X"88", X"0b", X"02", X"20", X"10", X"21", 
  X"8f", X"bf", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"3c", X"02", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"42", X"04", X"38", 
  X"3c", X"02", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8c", X"42", X"08", X"a0", X"3c", X"02", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"42", X"04", X"18", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"3c", X"02", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"24", X"42", X"04", X"58", X"3c", X"03", X"00", X"00", 
  X"00", X"80", X"10", X"21", X"8c", X"64", X"08", X"9c", 
  X"00", X"a0", X"30", X"21", X"0b", X"f0", X"0f", X"07", 
  X"00", X"40", X"28", X"21", X"3c", X"02", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"42", X"04", X"58", 
  X"94", X"a2", X"00", X"0c", X"27", X"bd", X"ff", X"98", 
  X"af", X"b0", X"00", X"54", X"30", X"42", X"00", X"02", 
  X"af", X"bf", X"00", X"64", X"af", X"b3", X"00", X"60", 
  X"af", X"b2", X"00", X"5c", X"af", X"b1", X"00", X"58", 
  X"14", X"40", X"00", X"2f", X"00", X"a0", X"80", X"21", 
  X"84", X"a5", X"00", X"0e", X"04", X"a1", X"00", X"0a", 
  X"00", X"80", X"90", X"21", X"86", X"02", X"00", X"0c", 
  X"24", X"11", X"00", X"40", X"24", X"03", X"04", X"00", 
  X"30", X"44", X"00", X"80", X"34", X"42", X"08", X"00", 
  X"00", X"64", X"88", X"0a", X"a6", X"02", X"00", X"0c", 
  X"0b", X"f0", X"0f", X"6b", X"00", X"00", X"98", X"21", 
  X"0f", X"f0", X"16", X"4b", X"27", X"a6", X"00", X"10", 
  X"04", X"40", X"ff", X"f4", X"8f", X"a3", X"00", X"14", 
  X"34", X"04", X"80", X"00", X"96", X"02", X"00", X"0c", 
  X"30", X"63", X"f0", X"00", X"38", X"73", X"20", X"00", 
  X"14", X"64", X"00", X"0b", X"2e", X"73", X"00", X"01", 
  X"8e", X"04", X"00", X"28", X"3c", X"03", X"bf", X"c0", 
  X"24", X"63", X"51", X"78", X"54", X"83", X"00", X"07", 
  X"34", X"42", X"08", X"00", X"34", X"42", X"04", X"00", 
  X"a6", X"02", X"00", X"0c", X"24", X"02", X"04", X"00", 
  X"0b", X"f0", X"0f", X"6a", X"ae", X"02", X"00", X"4c", 
  X"34", X"42", X"08", X"00", X"a6", X"02", X"00", X"0c", 
  X"24", X"11", X"04", X"00", X"02", X"40", X"20", X"21", 
  X"0f", X"f0", X"0f", X"94", X"02", X"20", X"28", X"21", 
  X"14", X"40", X"00", X"0d", X"3c", X"03", X"bf", X"c0", 
  X"86", X"02", X"00", X"0c", X"30", X"43", X"02", X"00", 
  X"14", X"60", X"00", X"1b", X"8f", X"bf", X"00", X"64", 
  X"34", X"42", X"00", X"02", X"a6", X"02", X"00", X"0c", 
  X"26", X"02", X"00", X"43", X"ae", X"02", X"00", X"00", 
  X"ae", X"02", X"00", X"10", X"24", X"02", X"00", X"01", 
  X"0b", X"f0", X"0f", X"8d", X"ae", X"02", X"00", X"14", 
  X"24", X"63", X"2d", X"ac", X"ae", X"43", X"00", X"3c", 
  X"96", X"03", X"00", X"0c", X"ae", X"02", X"00", X"00", 
  X"ae", X"02", X"00", X"10", X"34", X"63", X"00", X"80", 
  X"a6", X"03", X"00", X"0c", X"12", X"60", X"00", X"09", 
  X"ae", X"11", X"00", X"14", X"86", X"05", X"00", X"0e", 
  X"0f", X"f0", X"16", X"60", X"02", X"40", X"20", X"21", 
  X"10", X"40", X"00", X"05", X"8f", X"bf", X"00", X"64", 
  X"96", X"02", X"00", X"0c", X"34", X"42", X"00", X"01", 
  X"a6", X"02", X"00", X"0c", X"8f", X"bf", X"00", X"64", 
  X"8f", X"b3", X"00", X"60", X"8f", X"b2", X"00", X"5c", 
  X"8f", X"b1", X"00", X"58", X"8f", X"b0", X"00", X"54", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"68", 
  X"24", X"a2", X"00", X"0b", X"27", X"bd", X"ff", X"c0", 
  X"2c", X"43", X"00", X"17", X"af", X"b3", X"00", X"24", 
  X"af", X"bf", X"00", X"3c", X"af", X"be", X"00", X"38", 
  X"af", X"b7", X"00", X"34", X"af", X"b6", X"00", X"30", 
  X"af", X"b5", X"00", X"2c", X"af", X"b4", X"00", X"28", 
  X"af", X"b2", X"00", X"20", X"af", X"b1", X"00", X"1c", 
  X"af", X"b0", X"00", X"18", X"14", X"60", X"00", X"07", 
  X"00", X"80", X"98", X"21", X"24", X"11", X"ff", X"f8", 
  X"00", X"51", X"88", X"24", X"06", X"23", X"00", X"05", 
  X"02", X"25", X"28", X"2b", X"0b", X"f0", X"0f", X"ad", 
  X"24", X"02", X"00", X"0c", X"24", X"11", X"00", X"10", 
  X"02", X"25", X"28", X"2b", X"10", X"a0", X"00", X"03", 
  X"24", X"02", X"00", X"0c", X"0b", X"f0", X"11", X"2a", 
  X"ae", X"62", X"00", X"00", X"0f", X"f0", X"12", X"9e", 
  X"02", X"60", X"20", X"21", X"3c", X"10", X"00", X"00", 
  X"2e", X"22", X"01", X"f8", X"10", X"40", X"00", X"11", 
  X"26", X"10", X"04", X"90", X"02", X"11", X"10", X"21", 
  X"8c", X"52", X"00", X"0c", X"16", X"42", X"00", X"05", 
  X"00", X"11", X"28", X"c2", X"26", X"42", X"00", X"08", 
  X"8e", X"52", X"00", X"14", X"12", X"42", X"00", X"3a", 
  X"24", X"a5", X"00", X"02", X"8e", X"42", X"00", X"04", 
  X"24", X"03", X"ff", X"fc", X"8e", X"44", X"00", X"08", 
  X"00", X"62", X"10", X"24", X"8e", X"43", X"00", X"0c", 
  X"ac", X"83", X"00", X"0c", X"0b", X"f0", X"10", X"0f", 
  X"ac", X"64", X"00", X"08", X"00", X"11", X"12", X"42", 
  X"10", X"40", X"00", X"18", X"24", X"05", X"00", X"3f", 
  X"2c", X"43", X"00", X"05", X"10", X"60", X"00", X"04", 
  X"2c", X"43", X"00", X"15", X"00", X"11", X"29", X"82", 
  X"0b", X"f0", X"0f", X"df", X"24", X"a5", X"00", X"38", 
  X"14", X"60", X"00", X"10", X"24", X"45", X"00", X"5b", 
  X"2c", X"43", X"00", X"55", X"10", X"60", X"00", X"04", 
  X"2c", X"43", X"01", X"55", X"00", X"11", X"2b", X"02", 
  X"0b", X"f0", X"0f", X"df", X"24", X"a5", X"00", X"6e", 
  X"10", X"60", X"00", X"04", X"2c", X"42", X"05", X"55", 
  X"00", X"11", X"2b", X"c2", X"0b", X"f0", X"0f", X"df", 
  X"24", X"a5", X"00", X"77", X"10", X"40", X"00", X"03", 
  X"24", X"05", X"00", X"7e", X"00", X"11", X"2c", X"82", 
  X"24", X"a5", X"00", X"7c", X"00", X"05", X"10", X"c0", 
  X"02", X"02", X"10", X"21", X"8c", X"52", X"00", X"0c", 
  X"24", X"06", X"ff", X"fc", X"52", X"42", X"00", X"12", 
  X"24", X"a5", X"00", X"01", X"8e", X"43", X"00", X"04", 
  X"00", X"c3", X"18", X"24", X"00", X"71", X"20", X"23", 
  X"28", X"87", X"00", X"10", X"14", X"e0", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"0f", X"f5", 
  X"24", X"a5", X"ff", X"ff", X"04", X"82", X"ff", X"f5", 
  X"8e", X"52", X"00", X"0c", X"8e", X"42", X"00", X"0c", 
  X"8e", X"44", X"00", X"08", X"ac", X"82", X"00", X"0c", 
  X"ac", X"44", X"00", X"08", X"0b", X"f0", X"10", X"10", 
  X"02", X"43", X"10", X"21", X"24", X"a5", X"00", X"01", 
  X"8e", X"12", X"00", X"10", X"3c", X"04", X"00", X"00", 
  X"24", X"84", X"04", X"98", X"12", X"44", X"00", X"5a", 
  X"24", X"03", X"ff", X"fc", X"8e", X"42", X"00", X"04", 
  X"00", X"62", X"10", X"24", X"00", X"51", X"18", X"23", 
  X"28", X"66", X"00", X"10", X"54", X"c0", X"00", X"0d", 
  X"ae", X"04", X"00", X"14", X"02", X"51", X"10", X"21", 
  X"36", X"31", X"00", X"01", X"ae", X"51", X"00", X"04", 
  X"ae", X"02", X"00", X"14", X"ae", X"02", X"00", X"10", 
  X"ac", X"44", X"00", X"0c", X"ac", X"44", X"00", X"08", 
  X"34", X"64", X"00", X"01", X"ac", X"44", X"00", X"04", 
  X"00", X"43", X"10", X"21", X"0b", X"f0", X"11", X"32", 
  X"ac", X"43", X"00", X"00", X"04", X"60", X"00", X"06", 
  X"ae", X"04", X"00", X"10", X"02", X"42", X"10", X"21", 
  X"8c", X"43", X"00", X"04", X"34", X"63", X"00", X"01", 
  X"0b", X"f0", X"11", X"32", X"ac", X"43", X"00", X"04", 
  X"2c", X"43", X"02", X"00", X"10", X"60", X"00", X"0c", 
  X"00", X"02", X"32", X"42", X"00", X"02", X"10", X"c2", 
  X"00", X"02", X"18", X"83", X"24", X"06", X"00", X"01", 
  X"00", X"66", X"18", X"04", X"8e", X"06", X"00", X"04", 
  X"00", X"02", X"10", X"c0", X"02", X"02", X"10", X"21", 
  X"00", X"66", X"18", X"25", X"ae", X"03", X"00", X"04", 
  X"0b", X"f0", X"10", X"50", X"8c", X"43", X"00", X"08", 
  X"2c", X"c3", X"00", X"05", X"10", X"60", X"00", X"04", 
  X"2c", X"c3", X"00", X"15", X"00", X"02", X"31", X"82", 
  X"0b", X"f0", X"10", X"3a", X"24", X"c6", X"00", X"38", 
  X"10", X"60", X"00", X"03", X"2c", X"c3", X"00", X"55", 
  X"0b", X"f0", X"10", X"3a", X"24", X"c6", X"00", X"5b", 
  X"10", X"60", X"00", X"04", X"2c", X"c3", X"01", X"55", 
  X"00", X"02", X"33", X"02", X"0b", X"f0", X"10", X"3a", 
  X"24", X"c6", X"00", X"6e", X"10", X"60", X"00", X"04", 
  X"2c", X"c3", X"05", X"55", X"00", X"02", X"33", X"c2", 
  X"0b", X"f0", X"10", X"3a", X"24", X"c6", X"00", X"77", 
  X"10", X"60", X"00", X"03", X"24", X"06", X"00", X"7e", 
  X"00", X"02", X"34", X"82", X"24", X"c6", X"00", X"7c", 
  X"00", X"06", X"38", X"c0", X"02", X"07", X"38", X"21", 
  X"8c", X"e3", X"00", X"08", X"50", X"67", X"00", X"03", 
  X"24", X"02", X"00", X"01", X"0b", X"f0", X"10", X"4a", 
  X"24", X"08", X"ff", X"fc", X"00", X"06", X"30", X"83", 
  X"00", X"c2", X"30", X"04", X"8e", X"02", X"00", X"04", 
  X"00", X"c2", X"30", X"25", X"ae", X"06", X"00", X"04", 
  X"0b", X"f0", X"10", X"50", X"00", X"60", X"10", X"21", 
  X"50", X"67", X"00", X"07", X"8c", X"62", X"00", X"0c", 
  X"8c", X"66", X"00", X"04", X"01", X"06", X"30", X"24", 
  X"00", X"46", X"30", X"2b", X"54", X"c0", X"ff", X"fa", 
  X"8c", X"63", X"00", X"08", X"8c", X"62", X"00", X"0c", 
  X"ae", X"42", X"00", X"0c", X"ae", X"43", X"00", X"08", 
  X"ac", X"52", X"00", X"08", X"ac", X"72", X"00", X"0c", 
  X"00", X"05", X"10", X"83", X"24", X"03", X"00", X"01", 
  X"00", X"43", X"18", X"04", X"8e", X"02", X"00", X"04", 
  X"00", X"43", X"30", X"2b", X"54", X"c0", X"00", X"4f", 
  X"8e", X"14", X"00", X"08", X"00", X"62", X"30", X"24", 
  X"14", X"c0", X"00", X"08", X"24", X"0a", X"ff", X"fc", 
  X"24", X"06", X"ff", X"fc", X"00", X"a6", X"28", X"24", 
  X"00", X"03", X"18", X"40", X"00", X"62", X"30", X"24", 
  X"10", X"c0", X"ff", X"fd", X"24", X"a5", X"00", X"04", 
  X"24", X"0a", X"ff", X"fc", X"00", X"05", X"10", X"c0", 
  X"02", X"02", X"10", X"21", X"00", X"40", X"40", X"21", 
  X"00", X"a0", X"38", X"21", X"8d", X"12", X"00", X"0c", 
  X"52", X"48", X"00", X"22", X"24", X"e7", X"00", X"01", 
  X"8e", X"49", X"00", X"04", X"01", X"49", X"48", X"24", 
  X"01", X"31", X"30", X"23", X"28", X"cb", X"00", X"10", 
  X"15", X"60", X"00", X"11", X"00", X"00", X"00", X"00", 
  X"8e", X"43", X"00", X"0c", X"8e", X"45", X"00", X"08", 
  X"02", X"51", X"10", X"21", X"36", X"31", X"00", X"01", 
  X"ae", X"51", X"00", X"04", X"ac", X"a3", X"00", X"0c", 
  X"ac", X"65", X"00", X"08", X"34", X"c3", X"00", X"01", 
  X"ae", X"02", X"00", X"14", X"ae", X"02", X"00", X"10", 
  X"ac", X"44", X"00", X"0c", X"ac", X"44", X"00", X"08", 
  X"ac", X"43", X"00", X"04", X"00", X"46", X"10", X"21", 
  X"0b", X"f0", X"11", X"32", X"ac", X"46", X"00", X"00", 
  X"04", X"c2", X"ff", X"e7", X"8e", X"52", X"00", X"0c", 
  X"02", X"49", X"10", X"21", X"8c", X"43", X"00", X"04", 
  X"34", X"63", X"00", X"01", X"ac", X"43", X"00", X"04", 
  X"8e", X"42", X"00", X"0c", X"8e", X"43", X"00", X"08", 
  X"ac", X"62", X"00", X"0c", X"0b", X"f0", X"11", X"32", 
  X"ac", X"43", X"00", X"08", X"30", X"e6", X"00", X"03", 
  X"14", X"c0", X"ff", X"da", X"25", X"08", X"00", X"08", 
  X"30", X"a6", X"00", X"03", X"14", X"c0", X"00", X"06", 
  X"24", X"46", X"ff", X"f8", X"8e", X"05", X"00", X"04", 
  X"00", X"03", X"10", X"27", X"00", X"45", X"10", X"24", 
  X"0b", X"f0", X"10", X"9b", X"ae", X"02", X"00", X"04", 
  X"8c", X"42", X"00", X"00", X"10", X"46", X"ff", X"f6", 
  X"24", X"a5", X"ff", X"ff", X"8e", X"02", X"00", X"04", 
  X"00", X"03", X"18", X"40", X"00", X"43", X"28", X"2b", 
  X"54", X"a0", X"00", X"0a", X"8e", X"14", X"00", X"08", 
  X"10", X"60", X"00", X"07", X"00", X"e0", X"28", X"21", 
  X"00", X"62", X"30", X"24", X"54", X"c0", X"ff", X"c2", 
  X"00", X"05", X"10", X"c0", X"24", X"a5", X"00", X"04", 
  X"0b", X"f0", X"10", X"a2", X"00", X"03", X"18", X"40", 
  X"8e", X"14", X"00", X"08", X"24", X"15", X"ff", X"fc", 
  X"8e", X"82", X"00", X"04", X"02", X"a2", X"a8", X"24", 
  X"02", X"b1", X"10", X"2b", X"14", X"40", X"00", X"04", 
  X"02", X"b1", X"18", X"23", X"28", X"62", X"00", X"10", 
  X"50", X"40", X"00", X"7b", X"8e", X"12", X"00", X"08", 
  X"3c", X"02", X"00", X"00", X"8c", X"56", X"0d", X"5c", 
  X"3c", X"02", X"00", X"00", X"8c", X"44", X"08", X"a4", 
  X"00", X"40", X"18", X"21", X"24", X"02", X"ff", X"ff", 
  X"02", X"95", X"f0", X"21", X"14", X"82", X"00", X"03", 
  X"02", X"36", X"b0", X"21", X"0b", X"f0", X"10", X"c0", 
  X"26", X"d6", X"00", X"10", X"26", X"d6", X"10", X"0f", 
  X"24", X"02", X"f0", X"00", X"02", X"c2", X"b0", X"24", 
  X"02", X"60", X"20", X"21", X"02", X"c0", X"28", X"21", 
  X"0f", X"f0", X"14", X"15", X"af", X"a3", X"00", X"10", 
  X"00", X"40", X"90", X"21", X"24", X"02", X"ff", X"ff", 
  X"12", X"42", X"00", X"56", X"8f", X"a3", X"00", X"10", 
  X"02", X"5e", X"10", X"2b", X"10", X"40", X"00", X"04", 
  X"3c", X"17", X"00", X"00", X"56", X"90", X"00", X"52", 
  X"8e", X"02", X"00", X"08", X"3c", X"17", X"00", X"00", 
  X"8e", X"e2", X"08", X"cc", X"02", X"c2", X"10", X"21", 
  X"16", X"5e", X"00", X"09", X"ae", X"e2", X"08", X"cc", 
  X"32", X"44", X"0f", X"ff", X"14", X"80", X"00", X"07", 
  X"8c", X"64", X"08", X"a4", X"8e", X"02", X"00", X"08", 
  X"02", X"d5", X"a8", X"21", X"36", X"b5", X"00", X"01", 
  X"0b", X"f0", X"11", X"12", X"ac", X"55", X"00", X"04", 
  X"8c", X"64", X"08", X"a4", X"24", X"03", X"ff", X"ff", 
  X"54", X"83", X"00", X"04", X"02", X"5e", X"f0", X"23", 
  X"3c", X"02", X"00", X"00", X"0b", X"f0", X"10", X"e3", 
  X"ac", X"52", X"08", X"a4", X"00", X"5e", X"10", X"21", 
  X"ae", X"e2", X"08", X"cc", X"32", X"43", X"00", X"07", 
  X"10", X"60", X"00", X"04", X"00", X"00", X"10", X"21", 
  X"24", X"02", X"00", X"08", X"00", X"43", X"10", X"23", 
  X"02", X"42", X"90", X"21", X"02", X"56", X"b0", X"21", 
  X"24", X"42", X"10", X"00", X"32", X"d6", X"0f", X"ff", 
  X"00", X"56", X"b0", X"23", X"02", X"60", X"20", X"21", 
  X"0f", X"f0", X"14", X"15", X"02", X"c0", X"28", X"21", 
  X"24", X"03", X"ff", X"ff", X"14", X"43", X"00", X"03", 
  X"8e", X"e3", X"08", X"cc", X"02", X"40", X"10", X"21", 
  X"00", X"00", X"b0", X"21", X"00", X"52", X"10", X"23", 
  X"ae", X"12", X"00", X"08", X"02", X"c3", X"18", X"21", 
  X"00", X"56", X"b0", X"21", X"36", X"d6", X"00", X"01", 
  X"ae", X"e3", X"08", X"cc", X"12", X"90", X"00", X"16", 
  X"ae", X"56", X"00", X"04", X"2e", X"a2", X"00", X"10", 
  X"10", X"40", X"00", X"04", X"24", X"02", X"ff", X"f8", 
  X"24", X"02", X"00", X"01", X"0b", X"f0", X"11", X"1d", 
  X"ae", X"42", X"00", X"04", X"26", X"b5", X"ff", X"f4", 
  X"02", X"a2", X"a8", X"24", X"8e", X"82", X"00", X"04", 
  X"24", X"03", X"00", X"05", X"30", X"42", X"00", X"01", 
  X"02", X"a2", X"10", X"25", X"ae", X"82", X"00", X"04", 
  X"02", X"95", X"10", X"21", X"2e", X"b5", X"00", X"10", 
  X"ac", X"43", X"00", X"04", X"16", X"a0", X"00", X"04", 
  X"ac", X"43", X"00", X"08", X"02", X"60", X"20", X"21", 
  X"0f", X"f0", X"0c", X"ed", X"26", X"85", X"00", X"08", 
  X"3c", X"03", X"00", X"00", X"8e", X"e2", X"08", X"cc", 
  X"8c", X"64", X"0d", X"58", X"00", X"82", X"20", X"2b", 
  X"54", X"80", X"00", X"01", X"ac", X"62", X"0d", X"58", 
  X"3c", X"03", X"00", X"00", X"8c", X"64", X"0d", X"54", 
  X"00", X"82", X"20", X"2b", X"54", X"80", X"00", X"01", 
  X"ac", X"62", X"0d", X"54", X"8e", X"02", X"00", X"08", 
  X"24", X"03", X"ff", X"fc", X"8c", X"42", X"00", X"04", 
  X"00", X"62", X"10", X"24", X"00", X"51", X"18", X"23", 
  X"00", X"51", X"10", X"2b", X"14", X"40", X"00", X"04", 
  X"00", X"00", X"00", X"00", X"28", X"62", X"00", X"10", 
  X"50", X"40", X"00", X"05", X"8e", X"12", X"00", X"08", 
  X"0f", X"f0", X"12", X"a0", X"02", X"60", X"20", X"21", 
  X"0b", X"f0", X"11", X"35", X"00", X"00", X"10", X"21", 
  X"36", X"22", X"00", X"01", X"34", X"63", X"00", X"01", 
  X"02", X"51", X"88", X"21", X"ae", X"42", X"00", X"04", 
  X"ae", X"11", X"00", X"08", X"ae", X"23", X"00", X"04", 
  X"0f", X"f0", X"12", X"a0", X"02", X"60", X"20", X"21", 
  X"26", X"42", X"00", X"08", X"8f", X"bf", X"00", X"3c", 
  X"8f", X"be", X"00", X"38", X"8f", X"b7", X"00", X"34", 
  X"8f", X"b6", X"00", X"30", X"8f", X"b5", X"00", X"2c", 
  X"8f", X"b4", X"00", X"28", X"8f", X"b3", X"00", X"24", 
  X"8f", X"b2", X"00", X"20", X"8f", X"b1", X"00", X"1c", 
  X"8f", X"b0", X"00", X"18", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"40", X"30", X"a5", X"00", X"ff", 
  X"00", X"86", X"30", X"21", X"10", X"86", X"00", X"06", 
  X"00", X"00", X"00", X"00", X"90", X"82", X"00", X"00", 
  X"10", X"45", X"00", X"05", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"11", X"43", X"24", X"84", X"00", X"01", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"00", X"80", X"10", X"21", 
  X"28", X"ca", X"00", X"08", X"15", X"40", X"00", X"5f", 
  X"00", X"80", X"10", X"21", X"00", X"a4", X"c0", X"26", 
  X"33", X"18", X"00", X"03", X"17", X"00", X"00", X"64", 
  X"00", X"04", X"38", X"23", X"30", X"e7", X"00", X"03", 
  X"10", X"e0", X"00", X"05", X"00", X"c7", X"30", X"23", 
  X"88", X"b8", X"00", X"00", X"00", X"a7", X"28", X"21", 
  X"a8", X"98", X"00", X"00", X"00", X"87", X"20", X"21", 
  X"30", X"d8", X"00", X"3f", X"10", X"d8", X"00", X"32", 
  X"00", X"d8", X"38", X"23", X"00", X"87", X"38", X"21", 
  X"00", X"86", X"40", X"21", X"25", X"19", X"fe", X"e0", 
  X"cc", X"a4", X"00", X"00", X"cc", X"a4", X"00", X"20", 
  X"cc", X"a4", X"00", X"40", X"cc", X"a4", X"00", X"60", 
  X"8c", X"a8", X"00", X"00", X"03", X"24", X"18", X"2b", 
  X"1c", X"60", X"00", X"03", X"8c", X"a9", X"00", X"04", 
  X"cc", X"9e", X"00", X"80", X"cc", X"9e", X"00", X"a0", 
  X"8c", X"aa", X"00", X"08", X"8c", X"ab", X"00", X"0c", 
  X"8c", X"ac", X"00", X"10", X"8c", X"ad", X"00", X"14", 
  X"8c", X"ae", X"00", X"18", X"8c", X"af", X"00", X"1c", 
  X"cc", X"a4", X"00", X"80", X"ac", X"88", X"00", X"00", 
  X"ac", X"89", X"00", X"04", X"ac", X"8a", X"00", X"08", 
  X"ac", X"8b", X"00", X"0c", X"ac", X"8c", X"00", X"10", 
  X"ac", X"8d", X"00", X"14", X"ac", X"8e", X"00", X"18", 
  X"ac", X"8f", X"00", X"1c", X"8c", X"a8", X"00", X"20", 
  X"8c", X"a9", X"00", X"24", X"8c", X"aa", X"00", X"28", 
  X"8c", X"ab", X"00", X"2c", X"8c", X"ac", X"00", X"30", 
  X"8c", X"ad", X"00", X"34", X"8c", X"ae", X"00", X"38", 
  X"8c", X"af", X"00", X"3c", X"cc", X"a4", X"00", X"a0", 
  X"ac", X"88", X"00", X"20", X"ac", X"89", X"00", X"24", 
  X"ac", X"8a", X"00", X"28", X"ac", X"8b", X"00", X"2c", 
  X"ac", X"8c", X"00", X"30", X"ac", X"8d", X"00", X"34", 
  X"ac", X"8e", X"00", X"38", X"ac", X"8f", X"00", X"3c", 
  X"24", X"84", X"00", X"40", X"14", X"87", X"ff", X"d8", 
  X"24", X"a5", X"00", X"40", X"03", X"00", X"30", X"21", 
  X"cc", X"a4", X"00", X"00", X"30", X"d8", X"00", X"1f", 
  X"10", X"d8", X"00", X"13", X"00", X"00", X"00", X"00", 
  X"8c", X"a8", X"00", X"00", X"8c", X"a9", X"00", X"04", 
  X"8c", X"aa", X"00", X"08", X"8c", X"ab", X"00", X"0c", 
  X"8c", X"ac", X"00", X"10", X"8c", X"ad", X"00", X"14", 
  X"8c", X"ae", X"00", X"18", X"8c", X"af", X"00", X"1c", 
  X"24", X"a5", X"00", X"20", X"ac", X"88", X"00", X"00", 
  X"ac", X"89", X"00", X"04", X"ac", X"8a", X"00", X"08", 
  X"ac", X"8b", X"00", X"0c", X"ac", X"8c", X"00", X"10", 
  X"ac", X"8d", X"00", X"14", X"ac", X"8e", X"00", X"18", 
  X"ac", X"8f", X"00", X"1c", X"24", X"84", X"00", X"20", 
  X"33", X"06", X"00", X"03", X"10", X"d8", X"00", X"07", 
  X"03", X"06", X"38", X"23", X"00", X"87", X"38", X"21", 
  X"8c", X"ab", X"00", X"00", X"24", X"84", X"00", X"04", 
  X"24", X"a5", X"00", X"04", X"14", X"87", X"ff", X"fc", 
  X"ac", X"8b", X"ff", X"fc", X"18", X"c0", X"00", X"06", 
  X"00", X"86", X"38", X"21", X"80", X"a3", X"00", X"00", 
  X"24", X"84", X"00", X"01", X"24", X"a5", X"00", X"01", 
  X"14", X"87", X"ff", X"fc", X"a0", X"83", X"ff", X"ff", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"30", X"e7", X"00", X"03", X"10", X"e0", X"00", X"06", 
  X"00", X"c7", X"30", X"23", X"88", X"a3", X"00", X"00", 
  X"98", X"a3", X"00", X"03", X"00", X"a7", X"28", X"21", 
  X"a8", X"83", X"00", X"00", X"00", X"87", X"20", X"21", 
  X"30", X"d8", X"00", X"3f", X"10", X"d8", X"00", X"42", 
  X"00", X"d8", X"38", X"23", X"00", X"87", X"38", X"21", 
  X"00", X"86", X"40", X"21", X"25", X"19", X"fe", X"e0", 
  X"cc", X"a4", X"00", X"00", X"cc", X"a4", X"00", X"20", 
  X"cc", X"a4", X"00", X"40", X"cc", X"a4", X"00", X"60", 
  X"88", X"a8", X"00", X"00", X"88", X"a9", X"00", X"04", 
  X"88", X"aa", X"00", X"08", X"03", X"24", X"18", X"2b", 
  X"1c", X"60", X"00", X"03", X"88", X"ab", X"00", X"0c", 
  X"cc", X"9e", X"00", X"80", X"cc", X"9e", X"00", X"a0", 
  X"88", X"ac", X"00", X"10", X"88", X"ad", X"00", X"14", 
  X"88", X"ae", X"00", X"18", X"88", X"af", X"00", X"1c", 
  X"98", X"a8", X"00", X"03", X"98", X"a9", X"00", X"07", 
  X"98", X"aa", X"00", X"0b", X"98", X"ab", X"00", X"0f", 
  X"98", X"ac", X"00", X"13", X"98", X"ad", X"00", X"17", 
  X"98", X"ae", X"00", X"1b", X"98", X"af", X"00", X"1f", 
  X"cc", X"a4", X"00", X"80", X"ac", X"88", X"00", X"00", 
  X"ac", X"89", X"00", X"04", X"ac", X"8a", X"00", X"08", 
  X"ac", X"8b", X"00", X"0c", X"ac", X"8c", X"00", X"10", 
  X"ac", X"8d", X"00", X"14", X"ac", X"8e", X"00", X"18", 
  X"ac", X"8f", X"00", X"1c", X"88", X"a8", X"00", X"20", 
  X"88", X"a9", X"00", X"24", X"88", X"aa", X"00", X"28", 
  X"88", X"ab", X"00", X"2c", X"88", X"ac", X"00", X"30", 
  X"88", X"ad", X"00", X"34", X"88", X"ae", X"00", X"38", 
  X"88", X"af", X"00", X"3c", X"98", X"a8", X"00", X"23", 
  X"98", X"a9", X"00", X"27", X"98", X"aa", X"00", X"2b", 
  X"98", X"ab", X"00", X"2f", X"98", X"ac", X"00", X"33", 
  X"98", X"ad", X"00", X"37", X"98", X"ae", X"00", X"3b", 
  X"98", X"af", X"00", X"3f", X"cc", X"a4", X"00", X"a0", 
  X"ac", X"88", X"00", X"20", X"ac", X"89", X"00", X"24", 
  X"ac", X"8a", X"00", X"28", X"ac", X"8b", X"00", X"2c", 
  X"ac", X"8c", X"00", X"30", X"ac", X"8d", X"00", X"34", 
  X"ac", X"8e", X"00", X"38", X"ac", X"8f", X"00", X"3c", 
  X"24", X"84", X"00", X"40", X"14", X"87", X"ff", X"c7", 
  X"24", X"a5", X"00", X"40", X"03", X"00", X"30", X"21", 
  X"cc", X"a4", X"00", X"00", X"30", X"d8", X"00", X"1f", 
  X"10", X"d8", X"00", X"1b", X"00", X"00", X"00", X"00", 
  X"88", X"a8", X"00", X"00", X"88", X"a9", X"00", X"04", 
  X"88", X"aa", X"00", X"08", X"88", X"ab", X"00", X"0c", 
  X"88", X"ac", X"00", X"10", X"88", X"ad", X"00", X"14", 
  X"88", X"ae", X"00", X"18", X"88", X"af", X"00", X"1c", 
  X"98", X"a8", X"00", X"03", X"98", X"a9", X"00", X"07", 
  X"98", X"aa", X"00", X"0b", X"98", X"ab", X"00", X"0f", 
  X"98", X"ac", X"00", X"13", X"98", X"ad", X"00", X"17", 
  X"98", X"ae", X"00", X"1b", X"98", X"af", X"00", X"1f", 
  X"24", X"a5", X"00", X"20", X"ac", X"88", X"00", X"00", 
  X"ac", X"89", X"00", X"04", X"ac", X"8a", X"00", X"08", 
  X"ac", X"8b", X"00", X"0c", X"ac", X"8c", X"00", X"10", 
  X"ac", X"8d", X"00", X"14", X"ac", X"8e", X"00", X"18", 
  X"ac", X"8f", X"00", X"1c", X"24", X"84", X"00", X"20", 
  X"33", X"06", X"00", X"03", X"10", X"d8", X"00", X"08", 
  X"03", X"06", X"38", X"23", X"00", X"87", X"38", X"21", 
  X"88", X"a3", X"00", X"00", X"98", X"a3", X"00", X"03", 
  X"24", X"84", X"00", X"04", X"24", X"a5", X"00", X"04", 
  X"14", X"87", X"ff", X"fb", X"ac", X"83", X"ff", X"fc", 
  X"10", X"c0", X"ff", X"89", X"00", X"86", X"38", X"21", 
  X"80", X"a3", X"00", X"00", X"24", X"84", X"00", X"01", 
  X"24", X"a5", X"00", X"01", X"14", X"87", X"ff", X"fc", 
  X"a0", X"83", X"ff", X"ff", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"00", X"a4", X"18", X"2b", 
  X"14", X"60", X"00", X"03", X"00", X"80", X"10", X"21", 
  X"0b", X"f0", X"12", X"4a", X"00", X"00", X"18", X"21", 
  X"00", X"a6", X"20", X"21", X"00", X"44", X"18", X"2b", 
  X"10", X"60", X"00", X"0d", X"00", X"00", X"18", X"21", 
  X"00", X"06", X"18", X"23", X"00", X"46", X"38", X"21", 
  X"00", X"83", X"20", X"21", X"24", X"05", X"ff", X"ff", 
  X"00", X"e3", X"18", X"21", X"24", X"c6", X"ff", X"ff", 
  X"10", X"c5", X"00", X"0c", X"00", X"86", X"38", X"21", 
  X"90", X"e8", X"00", X"00", X"00", X"66", X"38", X"21", 
  X"0b", X"f0", X"12", X"43", X"a0", X"e8", X"00", X"00", 
  X"10", X"66", X"00", X"06", X"00", X"a3", X"20", X"21", 
  X"90", X"87", X"00", X"00", X"00", X"43", X"20", X"21", 
  X"24", X"63", X"00", X"01", X"0b", X"f0", X"12", X"4a", 
  X"a0", X"87", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"28", X"ca", X"00", X"08", 
  X"15", X"40", X"00", X"42", X"00", X"80", X"10", X"21", 
  X"10", X"a0", X"00", X"04", X"00", X"04", X"38", X"23", 
  X"00", X"00", X"00", X"00", X"7c", X"a5", X"7a", X"04", 
  X"7c", X"a5", X"fc", X"04", X"30", X"ea", X"00", X"03", 
  X"11", X"40", X"00", X"03", X"00", X"ca", X"30", X"23", 
  X"a8", X"85", X"00", X"00", X"00", X"8a", X"20", X"21", 
  X"30", X"ea", X"00", X"04", X"11", X"40", X"00", X"03", 
  X"00", X"ca", X"30", X"23", X"ac", X"85", X"00", X"00", 
  X"00", X"8a", X"20", X"21", X"30", X"d8", X"00", X"3f", 
  X"10", X"d8", X"00", X"1d", X"00", X"d8", X"38", X"23", 
  X"00", X"87", X"38", X"21", X"00", X"86", X"40", X"21", 
  X"25", X"19", X"fe", X"e0", X"03", X"24", X"18", X"2b", 
  X"1c", X"60", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"cc", X"9e", X"00", X"80", X"cc", X"9e", X"00", X"a0", 
  X"ac", X"85", X"00", X"00", X"ac", X"85", X"00", X"04", 
  X"ac", X"85", X"00", X"08", X"ac", X"85", X"00", X"0c", 
  X"ac", X"85", X"00", X"10", X"ac", X"85", X"00", X"14", 
  X"ac", X"85", X"00", X"18", X"ac", X"85", X"00", X"1c", 
  X"ac", X"85", X"00", X"20", X"ac", X"85", X"00", X"24", 
  X"ac", X"85", X"00", X"28", X"ac", X"85", X"00", X"2c", 
  X"ac", X"85", X"00", X"30", X"ac", X"85", X"00", X"34", 
  X"ac", X"85", X"00", X"38", X"ac", X"85", X"00", X"3c", 
  X"24", X"84", X"00", X"40", X"14", X"87", X"ff", X"e9", 
  X"00", X"00", X"00", X"00", X"03", X"00", X"30", X"21", 
  X"30", X"d8", X"00", X"1f", X"10", X"d8", X"00", X"0a", 
  X"00", X"00", X"00", X"00", X"ac", X"85", X"00", X"00", 
  X"ac", X"85", X"00", X"04", X"ac", X"85", X"00", X"08", 
  X"ac", X"85", X"00", X"0c", X"ac", X"85", X"00", X"10", 
  X"ac", X"85", X"00", X"14", X"ac", X"85", X"00", X"18", 
  X"ac", X"85", X"00", X"1c", X"24", X"84", X"00", X"20", 
  X"33", X"06", X"00", X"03", X"10", X"d8", X"00", X"05", 
  X"03", X"06", X"38", X"23", X"00", X"87", X"38", X"21", 
  X"24", X"84", X"00", X"04", X"14", X"87", X"ff", X"fe", 
  X"ac", X"85", X"ff", X"fc", X"18", X"c0", X"00", X"04", 
  X"00", X"86", X"38", X"21", X"24", X"84", X"00", X"01", 
  X"14", X"87", X"ff", X"fe", X"a0", X"85", X"ff", X"ff", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"27", X"bd", X"ff", X"c0", X"af", X"b0", X"00", X"18", 
  X"00", X"a0", X"80", X"21", X"af", X"bf", X"00", X"3c", 
  X"af", X"be", X"00", X"38", X"af", X"b7", X"00", X"34", 
  X"af", X"b6", X"00", X"30", X"af", X"b5", X"00", X"2c", 
  X"af", X"b4", X"00", X"28", X"af", X"b3", X"00", X"24", 
  X"af", X"b2", X"00", X"20", X"af", X"b1", X"00", X"1c", 
  X"16", X"00", X"00", X"05", X"00", X"c0", X"28", X"21", 
  X"0f", X"f0", X"0f", X"94", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"14", X"0a", X"8f", X"bf", X"00", X"3c", 
  X"00", X"80", X"a8", X"21", X"0f", X"f0", X"12", X"9e", 
  X"af", X"a6", X"00", X"10", X"8f", X"a5", X"00", X"10", 
  X"8e", X"07", X"ff", X"fc", X"24", X"13", X"ff", X"fc", 
  X"24", X"a2", X"00", X"0b", X"2c", X"43", X"00", X"17", 
  X"26", X"14", X"ff", X"f8", X"14", X"60", X"00", X"07", 
  X"00", X"f3", X"98", X"24", X"24", X"12", X"ff", X"f8", 
  X"00", X"52", X"90", X"24", X"06", X"43", X"00", X"05", 
  X"02", X"45", X"10", X"2b", X"0b", X"f0", X"12", X"ca", 
  X"24", X"02", X"00", X"0c", X"24", X"12", X"00", X"10", 
  X"02", X"45", X"10", X"2b", X"50", X"40", X"00", X"04", 
  X"02", X"72", X"10", X"2a", X"24", X"02", X"00", X"0c", 
  X"0b", X"f0", X"13", X"ae", X"ae", X"a2", X"00", X"00", 
  X"10", X"40", X"01", X"20", X"02", X"72", X"10", X"23", 
  X"3c", X"1e", X"00", X"00", X"27", X"de", X"04", X"90", 
  X"8f", X"c6", X"00", X"08", X"02", X"93", X"10", X"21", 
  X"10", X"46", X"00", X"08", X"8c", X"43", X"00", X"04", 
  X"24", X"04", X"ff", X"fe", X"00", X"83", X"20", X"24", 
  X"00", X"44", X"20", X"21", X"8c", X"84", X"00", X"04", 
  X"30", X"84", X"00", X"01", X"54", X"80", X"00", X"1f", 
  X"00", X"00", X"18", X"21", X"24", X"04", X"ff", X"fc", 
  X"00", X"83", X"18", X"24", X"14", X"46", X"00", X"12", 
  X"00", X"73", X"20", X"21", X"26", X"48", X"00", X"10", 
  X"00", X"88", X"40", X"2a", X"15", X"00", X"00", X"19", 
  X"30", X"e7", X"00", X"01", X"00", X"92", X"20", X"23", 
  X"02", X"92", X"a0", X"21", X"34", X"84", X"00", X"01", 
  X"af", X"d4", X"00", X"08", X"ae", X"84", X"00", X"04", 
  X"8e", X"02", X"ff", X"fc", X"02", X"a0", X"20", X"21", 
  X"30", X"42", X"00", X"01", X"02", X"42", X"90", X"25", 
  X"0f", X"f0", X"12", X"a0", X"ae", X"12", X"ff", X"fc", 
  X"0b", X"f0", X"14", X"09", X"02", X"00", X"10", X"21", 
  X"00", X"92", X"40", X"2a", X"15", X"00", X"00", X"09", 
  X"30", X"e7", X"00", X"01", X"8c", X"43", X"00", X"0c", 
  X"8c", X"42", X"00", X"08", X"00", X"80", X"98", X"21", 
  X"ac", X"43", X"00", X"0c", X"0b", X"f0", X"13", X"ec", 
  X"ac", X"62", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"30", X"e7", X"00", X"01", X"14", X"e0", X"00", X"ac", 
  X"24", X"16", X"ff", X"fc", X"8e", X"11", X"ff", X"f8", 
  X"02", X"91", X"88", X"23", X"8e", X"24", X"00", X"04", 
  X"02", X"c4", X"b0", X"24", X"10", X"40", X"00", X"75", 
  X"02", X"d3", X"b0", X"21", X"14", X"46", X"00", X"3f", 
  X"02", X"c3", X"b8", X"21", X"26", X"42", X"00", X"10", 
  X"02", X"e2", X"10", X"2a", X"14", X"40", X"00", X"70", 
  X"02", X"d2", X"10", X"2a", X"8e", X"22", X"00", X"0c", 
  X"8e", X"23", X"00", X"08", X"26", X"66", X"ff", X"fc", 
  X"ac", X"62", X"00", X"0c", X"ac", X"43", X"00", X"08", 
  X"2c", X"c2", X"00", X"25", X"10", X"40", X"00", X"23", 
  X"26", X"34", X"00", X"08", X"2c", X"c2", X"00", X"14", 
  X"14", X"40", X"00", X"19", X"02", X"80", X"18", X"21", 
  X"8e", X"02", X"00", X"00", X"ae", X"22", X"00", X"08", 
  X"8e", X"02", X"00", X"04", X"ae", X"22", X"00", X"0c", 
  X"2c", X"c2", X"00", X"1c", X"50", X"40", X"00", X"04", 
  X"8e", X"02", X"00", X"08", X"26", X"23", X"00", X"10", 
  X"0b", X"f0", X"13", X"2c", X"26", X"10", X"00", X"08", 
  X"ae", X"22", X"00", X"10", X"8e", X"02", X"00", X"0c", 
  X"ae", X"22", X"00", X"14", X"24", X"02", X"00", X"24", 
  X"50", X"c2", X"00", X"04", X"8e", X"02", X"00", X"10", 
  X"26", X"23", X"00", X"18", X"0b", X"f0", X"13", X"2c", 
  X"26", X"10", X"00", X"10", X"26", X"23", X"00", X"20", 
  X"26", X"10", X"00", X"18", X"ae", X"22", X"00", X"18", 
  X"8e", X"02", X"ff", X"fc", X"ae", X"22", X"00", X"1c", 
  X"8e", X"02", X"00", X"00", X"ac", X"62", X"00", X"00", 
  X"8e", X"02", X"00", X"04", X"ac", X"62", X"00", X"04", 
  X"8e", X"02", X"00", X"08", X"0b", X"f0", X"13", X"36", 
  X"ac", X"62", X"00", X"08", X"02", X"80", X"20", X"21", 
  X"0f", X"f0", X"12", X"35", X"02", X"00", X"28", X"21", 
  X"02", X"f2", X"b8", X"23", X"02", X"32", X"10", X"21", 
  X"36", X"f7", X"00", X"01", X"af", X"c2", X"00", X"08", 
  X"ac", X"57", X"00", X"04", X"8e", X"22", X"00", X"04", 
  X"02", X"a0", X"20", X"21", X"30", X"42", X"00", X"01", 
  X"02", X"42", X"90", X"25", X"0f", X"f0", X"12", X"a0", 
  X"ae", X"32", X"00", X"04", X"0b", X"f0", X"14", X"09", 
  X"02", X"80", X"10", X"21", X"02", X"f2", X"18", X"2a", 
  X"54", X"60", X"00", X"33", X"02", X"d2", X"10", X"2a", 
  X"8c", X"43", X"00", X"0c", X"8c", X"42", X"00", X"08", 
  X"26", X"66", X"ff", X"fc", X"ac", X"43", X"00", X"0c", 
  X"ac", X"62", X"00", X"08", X"8e", X"23", X"00", X"08", 
  X"8e", X"22", X"00", X"0c", X"ac", X"62", X"00", X"0c", 
  X"ac", X"43", X"00", X"08", X"2c", X"c2", X"00", X"25", 
  X"10", X"40", X"00", X"22", X"26", X"24", X"00", X"08", 
  X"2c", X"c2", X"00", X"14", X"14", X"40", X"00", X"19", 
  X"8e", X"02", X"00", X"00", X"ae", X"22", X"00", X"08", 
  X"8e", X"02", X"00", X"04", X"ae", X"22", X"00", X"0c", 
  X"2c", X"c2", X"00", X"1c", X"50", X"40", X"00", X"04", 
  X"8e", X"02", X"00", X"08", X"26", X"24", X"00", X"10", 
  X"0b", X"f0", X"13", X"6c", X"26", X"10", X"00", X"08", 
  X"ae", X"22", X"00", X"10", X"8e", X"02", X"00", X"0c", 
  X"ae", X"22", X"00", X"14", X"24", X"02", X"00", X"24", 
  X"50", X"c2", X"00", X"04", X"8e", X"02", X"00", X"10", 
  X"26", X"24", X"00", X"18", X"0b", X"f0", X"13", X"6c", 
  X"26", X"10", X"00", X"10", X"26", X"24", X"00", X"20", 
  X"26", X"10", X"00", X"18", X"ae", X"22", X"00", X"18", 
  X"8e", X"02", X"ff", X"fc", X"ae", X"22", X"00", X"1c", 
  X"8e", X"02", X"00", X"00", X"ac", X"82", X"00", X"00", 
  X"8e", X"02", X"00", X"04", X"ac", X"82", X"00", X"04", 
  X"8e", X"02", X"00", X"08", X"0b", X"f0", X"13", X"75", 
  X"ac", X"82", X"00", X"08", X"0f", X"f0", X"12", X"35", 
  X"02", X"00", X"28", X"21", X"0b", X"f0", X"13", X"a2", 
  X"02", X"e0", X"98", X"21", X"02", X"d2", X"10", X"2a", 
  X"14", X"40", X"00", X"2f", X"26", X"66", X"ff", X"fc", 
  X"8e", X"22", X"00", X"0c", X"8e", X"23", X"00", X"08", 
  X"ac", X"62", X"00", X"0c", X"ac", X"43", X"00", X"08", 
  X"2c", X"c2", X"00", X"25", X"10", X"40", X"00", X"24", 
  X"26", X"24", X"00", X"08", X"2c", X"c2", X"00", X"14", 
  X"14", X"40", X"00", X"19", X"8e", X"02", X"00", X"00", 
  X"ae", X"22", X"00", X"08", X"8e", X"02", X"00", X"04", 
  X"ae", X"22", X"00", X"0c", X"2c", X"c2", X"00", X"1c", 
  X"50", X"40", X"00", X"04", X"8e", X"02", X"00", X"08", 
  X"26", X"24", X"00", X"10", X"0b", X"f0", X"13", X"9b", 
  X"26", X"10", X"00", X"08", X"ae", X"22", X"00", X"10", 
  X"8e", X"02", X"00", X"0c", X"ae", X"22", X"00", X"14", 
  X"24", X"02", X"00", X"24", X"50", X"c2", X"00", X"04", 
  X"8e", X"02", X"00", X"10", X"26", X"24", X"00", X"18", 
  X"0b", X"f0", X"13", X"9b", X"26", X"10", X"00", X"10", 
  X"26", X"24", X"00", X"20", X"26", X"10", X"00", X"18", 
  X"ae", X"22", X"00", X"18", X"8e", X"02", X"ff", X"fc", 
  X"ae", X"22", X"00", X"1c", X"8e", X"02", X"00", X"00", 
  X"ac", X"82", X"00", X"00", X"8e", X"02", X"00", X"04", 
  X"ac", X"82", X"00", X"04", X"8e", X"02", X"00", X"08", 
  X"ac", X"82", X"00", X"08", X"02", X"c0", X"98", X"21", 
  X"0b", X"f0", X"13", X"ec", X"02", X"20", X"a0", X"21", 
  X"0f", X"f0", X"12", X"35", X"02", X"00", X"28", X"21", 
  X"0b", X"f0", X"13", X"a2", X"02", X"c0", X"98", X"21", 
  X"0f", X"f0", X"0f", X"94", X"02", X"a0", X"20", X"21", 
  X"14", X"40", X"00", X"05", X"00", X"40", X"88", X"21", 
  X"0f", X"f0", X"12", X"a0", X"02", X"a0", X"20", X"21", 
  X"0b", X"f0", X"14", X"09", X"00", X"00", X"10", X"21", 
  X"24", X"43", X"ff", X"f8", X"8e", X"02", X"ff", X"fc", 
  X"24", X"04", X"ff", X"fe", X"00", X"82", X"10", X"24", 
  X"02", X"82", X"10", X"21", X"14", X"62", X"00", X"06", 
  X"26", X"66", X"ff", X"fc", X"8e", X"22", X"ff", X"fc", 
  X"24", X"03", X"ff", X"fc", X"00", X"62", X"10", X"24", 
  X"0b", X"f0", X"13", X"ec", X"02", X"62", X"98", X"21", 
  X"2c", X"c2", X"00", X"25", X"10", X"40", X"00", X"25", 
  X"02", X"20", X"20", X"21", X"2c", X"c2", X"00", X"14", 
  X"14", X"40", X"00", X"1a", X"02", X"20", X"10", X"21", 
  X"8e", X"02", X"00", X"00", X"ae", X"22", X"00", X"00", 
  X"8e", X"02", X"00", X"04", X"ae", X"22", X"00", X"04", 
  X"2c", X"c2", X"00", X"1c", X"50", X"40", X"00", X"04", 
  X"8e", X"02", X"00", X"08", X"26", X"22", X"00", X"08", 
  X"0b", X"f0", X"13", X"dc", X"26", X"03", X"00", X"08", 
  X"ae", X"22", X"00", X"08", X"8e", X"02", X"00", X"0c", 
  X"ae", X"22", X"00", X"0c", X"24", X"02", X"00", X"24", 
  X"50", X"c2", X"00", X"04", X"8e", X"02", X"00", X"10", 
  X"26", X"22", X"00", X"10", X"0b", X"f0", X"13", X"dc", 
  X"26", X"03", X"00", X"10", X"26", X"03", X"00", X"18", 
  X"ae", X"22", X"00", X"10", X"8e", X"04", X"00", X"14", 
  X"26", X"22", X"00", X"18", X"0b", X"f0", X"13", X"dc", 
  X"ae", X"24", X"00", X"14", X"02", X"00", X"18", X"21", 
  X"8c", X"64", X"00", X"00", X"ac", X"44", X"00", X"00", 
  X"8c", X"64", X"00", X"04", X"ac", X"44", X"00", X"04", 
  X"8c", X"63", X"00", X"08", X"0b", X"f0", X"13", X"e5", 
  X"ac", X"43", X"00", X"08", X"0f", X"f0", X"12", X"35", 
  X"02", X"00", X"28", X"21", X"02", X"a0", X"20", X"21", 
  X"0f", X"f0", X"0c", X"ed", X"02", X"00", X"28", X"21", 
  X"0f", X"f0", X"12", X"a0", X"02", X"a0", X"20", X"21", 
  X"0b", X"f0", X"14", X"09", X"02", X"20", X"10", X"21", 
  X"02", X"72", X"10", X"23", X"2c", X"44", X"00", X"10", 
  X"14", X"80", X"00", X"10", X"8e", X"83", X"00", X"04", 
  X"30", X"63", X"00", X"01", X"02", X"92", X"28", X"21", 
  X"02", X"43", X"90", X"25", X"34", X"43", X"00", X"01", 
  X"ae", X"92", X"00", X"04", X"00", X"a2", X"10", X"21", 
  X"ac", X"a3", X"00", X"04", X"8c", X"43", X"00", X"04", 
  X"02", X"a0", X"20", X"21", X"24", X"a5", X"00", X"08", 
  X"34", X"63", X"00", X"01", X"0f", X"f0", X"0c", X"ed", 
  X"ac", X"43", X"00", X"04", X"0b", X"f0", X"14", X"06", 
  X"00", X"00", X"00", X"00", X"30", X"63", X"00", X"01", 
  X"02", X"63", X"18", X"25", X"ae", X"83", X"00", X"04", 
  X"02", X"93", X"98", X"21", X"8e", X"62", X"00", X"04", 
  X"34", X"42", X"00", X"01", X"ae", X"62", X"00", X"04", 
  X"0f", X"f0", X"12", X"a0", X"02", X"a0", X"20", X"21", 
  X"26", X"82", X"00", X"08", X"8f", X"bf", X"00", X"3c", 
  X"8f", X"be", X"00", X"38", X"8f", X"b7", X"00", X"34", 
  X"8f", X"b6", X"00", X"30", X"8f", X"b5", X"00", X"2c", 
  X"8f", X"b4", X"00", X"28", X"8f", X"b3", X"00", X"24", 
  X"8f", X"b2", X"00", X"20", X"8f", X"b1", X"00", X"1c", 
  X"8f", X"b0", X"00", X"18", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"40", X"27", X"bd", X"ff", X"e0", 
  X"af", X"b1", X"00", X"18", X"af", X"b0", X"00", X"14", 
  X"00", X"80", X"88", X"21", X"3c", X"10", X"00", X"00", 
  X"00", X"a0", X"20", X"21", X"af", X"bf", X"00", X"1c", 
  X"0f", X"f0", X"06", X"45", X"ae", X"00", X"0d", X"44", 
  X"24", X"03", X"ff", X"ff", X"14", X"43", X"00", X"05", 
  X"8f", X"bf", X"00", X"1c", X"8e", X"03", X"0d", X"44", 
  X"54", X"60", X"00", X"01", X"ae", X"23", X"00", X"00", 
  X"8f", X"bf", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"27", X"bd", X"ff", X"e8", 
  X"af", X"b0", X"00", X"10", X"00", X"a0", X"80", X"21", 
  X"84", X"a5", X"00", X"0e", X"af", X"bf", X"00", X"14", 
  X"0f", X"f0", X"16", X"8a", X"00", X"00", X"00", X"00", 
  X"04", X"42", X"00", X"05", X"96", X"03", X"00", X"0c", 
  X"8e", X"03", X"00", X"50", X"00", X"62", X"18", X"21", 
  X"0b", X"f0", X"14", X"38", X"ae", X"03", X"00", X"50", 
  X"30", X"63", X"ef", X"ff", X"a6", X"03", X"00", X"0c", 
  X"8f", X"bf", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"18", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"94", X"a2", X"00", X"0c", X"27", X"bd", X"ff", X"d8", 
  X"af", X"b3", X"00", X"20", X"30", X"42", X"01", X"00", 
  X"af", X"b2", X"00", X"1c", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"af", X"bf", X"00", X"24", 
  X"00", X"80", X"98", X"21", X"00", X"a0", X"80", X"21", 
  X"00", X"c0", X"90", X"21", X"10", X"40", X"00", X"05", 
  X"00", X"e0", X"88", X"21", X"84", X"a5", X"00", X"0e", 
  X"00", X"00", X"30", X"21", X"0f", X"f0", X"16", X"74", 
  X"24", X"07", X"00", X"02", X"96", X"02", X"00", X"0c", 
  X"86", X"05", X"00", X"0e", X"02", X"60", X"20", X"21", 
  X"30", X"42", X"ef", X"ff", X"a6", X"02", X"00", X"0c", 
  X"02", X"40", X"30", X"21", X"0f", X"f0", X"15", X"e0", 
  X"02", X"20", X"38", X"21", X"8f", X"bf", X"00", X"24", 
  X"8f", X"b3", X"00", X"20", X"8f", X"b2", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"27", X"bd", X"ff", X"e8", X"af", X"b0", X"00", X"10", 
  X"00", X"a0", X"80", X"21", X"84", X"a5", X"00", X"0e", 
  X"af", X"bf", X"00", X"14", X"0f", X"f0", X"16", X"74", 
  X"00", X"00", X"00", X"00", X"24", X"04", X"ff", X"ff", 
  X"14", X"44", X"00", X"04", X"96", X"03", X"00", X"0c", 
  X"30", X"63", X"ef", X"ff", X"0b", X"f0", X"14", X"6e", 
  X"a6", X"03", X"00", X"0c", X"34", X"63", X"10", X"00", 
  X"a6", X"03", X"00", X"0c", X"ae", X"02", X"00", X"50", 
  X"8f", X"bf", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"18", 
  X"84", X"a5", X"00", X"0e", X"27", X"bd", X"ff", X"e8", 
  X"af", X"bf", X"00", X"14", X"0f", X"f0", X"15", X"f6", 
  X"00", X"00", X"00", X"00", X"8f", X"bf", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"18", 
  X"00", X"85", X"40", X"25", X"3c", X"09", X"01", X"01", 
  X"31", X"08", X"00", X"03", X"3c", X"0f", X"7f", X"7f", 
  X"15", X"00", X"00", X"56", X"35", X"29", X"01", X"01", 
  X"35", X"ef", X"7f", X"7f", X"8c", X"82", X"00", X"00", 
  X"8c", X"a3", X"00", X"00", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"3e", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"3a", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"04", 
  X"8c", X"a3", X"00", X"04", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"36", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"32", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"08", 
  X"8c", X"a3", X"00", X"08", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"2e", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"2a", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"0c", 
  X"8c", X"a3", X"00", X"0c", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"26", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"22", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"10", 
  X"8c", X"a3", X"00", X"10", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"1e", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"1a", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"14", 
  X"8c", X"a3", X"00", X"14", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"16", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"12", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"18", 
  X"8c", X"a3", X"00", X"18", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"0e", 
  X"01", X"0a", X"40", X"24", X"15", X"00", X"00", X"0a", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"1c", 
  X"8c", X"a3", X"00", X"1c", X"00", X"49", X"40", X"23", 
  X"00", X"4f", X"50", X"27", X"14", X"43", X"00", X"06", 
  X"01", X"0a", X"40", X"24", X"24", X"84", X"00", X"20", 
  X"11", X"00", X"ff", X"c0", X"24", X"a5", X"00", X"20", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"00", X"43", X"50", X"26", X"01", X"48", X"58", X"25", 
  X"00", X"0b", X"74", X"02", X"15", X"c0", X"00", X"04", 
  X"00", X"00", X"00", X"00", X"00", X"0b", X"5c", X"00", 
  X"00", X"02", X"14", X"00", X"00", X"03", X"1c", X"00", 
  X"00", X"0b", X"76", X"02", X"15", X"c0", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"00", X"02", X"12", X"00", 
  X"00", X"03", X"1a", X"00", X"00", X"02", X"16", X"02", 
  X"00", X"03", X"1e", X"02", X"03", X"e0", X"00", X"08", 
  X"00", X"43", X"10", X"23", X"90", X"88", X"00", X"00", 
  X"90", X"a9", X"00", X"00", X"11", X"00", X"00", X"03", 
  X"24", X"84", X"00", X"01", X"11", X"09", X"ff", X"fb", 
  X"24", X"a5", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"01", X"09", X"10", X"23", X"90", X"8a", X"00", X"00", 
  X"00", X"80", X"10", X"21", X"15", X"40", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"24", X"02", X"00", X"00", X"90", X"8a", X"00", X"01", 
  X"15", X"40", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"00", X"01", 
  X"90", X"8a", X"00", X"02", X"15", X"40", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"24", X"02", X"00", X"02", X"90", X"8a", X"00", X"03", 
  X"15", X"40", X"00", X"03", X"00", X"04", X"20", X"82", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"00", X"03", 
  X"24", X"84", X"00", X"01", X"00", X"04", X"20", X"80", 
  X"8c", X"8a", X"00", X"00", X"3c", X"09", X"01", X"01", 
  X"35", X"29", X"01", X"01", X"00", X"09", X"79", X"c0", 
  X"01", X"49", X"40", X"23", X"01", X"0f", X"40", X"24", 
  X"11", X"00", X"00", X"06", X"01", X"0a", X"60", X"24", 
  X"11", X"88", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"90", X"8a", X"00", X"00", X"10", X"00", X"00", X"22", 
  X"24", X"84", X"00", X"00", X"8c", X"8b", X"00", X"04", 
  X"01", X"69", X"40", X"23", X"01", X"0f", X"40", X"24", 
  X"11", X"00", X"00", X"06", X"01", X"0b", X"60", X"24", 
  X"11", X"88", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"90", X"8a", X"00", X"04", X"10", X"00", X"00", X"18", 
  X"24", X"84", X"00", X"04", X"8c", X"8a", X"00", X"08", 
  X"01", X"49", X"40", X"23", X"01", X"0f", X"40", X"24", 
  X"11", X"00", X"00", X"06", X"01", X"0a", X"60", X"24", 
  X"11", X"88", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"90", X"8a", X"00", X"08", X"10", X"00", X"00", X"0e", 
  X"24", X"84", X"00", X"08", X"8c", X"8b", X"00", X"0c", 
  X"01", X"69", X"40", X"23", X"01", X"0f", X"40", X"24", 
  X"11", X"00", X"00", X"06", X"01", X"0b", X"60", X"24", 
  X"11", X"88", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"90", X"8a", X"00", X"0c", X"10", X"00", X"00", X"04", 
  X"24", X"84", X"00", X"0c", X"8c", X"8a", X"00", X"10", 
  X"10", X"00", X"ff", X"d7", X"24", X"84", X"00", X"10", 
  X"15", X"40", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"24", X"84", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"82", X"10", X"23", X"90", X"8a", X"00", X"01", 
  X"15", X"40", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"24", X"84", X"00", X"01", X"03", X"e0", X"00", X"08", 
  X"00", X"82", X"10", X"23", X"90", X"8a", X"00", X"02", 
  X"15", X"40", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"24", X"84", X"00", X"02", X"03", X"e0", X"00", X"08", 
  X"00", X"82", X"10", X"23", X"90", X"8a", X"00", X"03", 
  X"24", X"84", X"00", X"03", X"03", X"e0", X"00", X"08", 
  X"00", X"82", X"10", X"23", X"27", X"bd", X"ff", X"e0", 
  X"af", X"b2", X"00", X"18", X"af", X"b1", X"00", X"14", 
  X"af", X"b0", X"00", X"10", X"af", X"bf", X"00", X"1c", 
  X"00", X"80", X"88", X"21", X"00", X"a0", X"90", X"21", 
  X"10", X"80", X"00", X"06", X"00", X"c0", X"80", X"21", 
  X"8c", X"82", X"00", X"38", X"54", X"40", X"00", X"04", 
  X"8e", X"02", X"00", X"18", X"0f", X"f0", X"0b", X"91", 
  X"00", X"00", X"00", X"00", X"8e", X"02", X"00", X"18", 
  X"ae", X"02", X"00", X"08", X"96", X"02", X"00", X"0c", 
  X"30", X"42", X"00", X"08", X"10", X"40", X"00", X"0f", 
  X"02", X"20", X"20", X"21", X"8e", X"02", X"00", X"10", 
  X"10", X"40", X"00", X"0c", X"00", X"00", X"00", X"00", 
  X"86", X"02", X"00", X"0c", X"30", X"43", X"20", X"00", 
  X"14", X"60", X"00", X"0e", X"32", X"52", X"00", X"ff", 
  X"8e", X"03", X"00", X"60", X"34", X"42", X"20", X"00", 
  X"a6", X"02", X"00", X"0c", X"24", X"02", X"df", X"ff", 
  X"00", X"62", X"10", X"24", X"0b", X"f0", X"15", X"5f", 
  X"ae", X"02", X"00", X"60", X"0f", X"f0", X"0a", X"69", 
  X"02", X"00", X"28", X"21", X"50", X"40", X"ff", X"f3", 
  X"86", X"02", X"00", X"0c", X"0b", X"f0", X"15", X"83", 
  X"24", X"02", X"ff", X"ff", X"8e", X"03", X"00", X"00", 
  X"8e", X"02", X"00", X"10", X"00", X"62", X"10", X"23", 
  X"8e", X"03", X"00", X"14", X"00", X"43", X"18", X"2a", 
  X"54", X"60", X"00", X"07", X"8e", X"03", X"00", X"08", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"0b", X"46", 
  X"02", X"00", X"28", X"21", X"54", X"40", X"00", X"19", 
  X"24", X"02", X"ff", X"ff", X"8e", X"03", X"00", X"08", 
  X"24", X"42", X"00", X"01", X"24", X"63", X"ff", X"ff", 
  X"ae", X"03", X"00", X"08", X"8e", X"03", X"00", X"00", 
  X"24", X"64", X"00", X"01", X"ae", X"04", X"00", X"00", 
  X"a0", X"72", X"00", X"00", X"8e", X"03", X"00", X"14", 
  X"50", X"43", X"00", X"09", X"02", X"20", X"20", X"21", 
  X"96", X"03", X"00", X"0c", X"30", X"63", X"00", X"01", 
  X"10", X"60", X"00", X"0a", X"02", X"40", X"10", X"21", 
  X"24", X"03", X"00", X"0a", X"16", X"43", X"00", X"08", 
  X"8f", X"bf", X"00", X"1c", X"02", X"20", X"20", X"21", 
  X"0f", X"f0", X"0b", X"46", X"02", X"00", X"28", X"21", 
  X"14", X"40", X"00", X"02", X"24", X"02", X"ff", X"ff", 
  X"02", X"40", X"10", X"21", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b2", X"00", X"18", X"8f", X"b1", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"3c", X"03", X"00", X"00", 
  X"00", X"80", X"10", X"21", X"8c", X"64", X"08", X"9c", 
  X"00", X"a0", X"30", X"21", X"0b", X"f0", X"15", X"37", 
  X"00", X"40", X"28", X"21", X"27", X"bd", X"ff", X"c0", 
  X"3c", X"02", X"00", X"00", X"af", X"b2", X"00", X"38", 
  X"af", X"b1", X"00", X"34", X"af", X"b0", X"00", X"30", 
  X"af", X"bf", X"00", X"3c", X"00", X"80", X"80", X"21", 
  X"00", X"e0", X"88", X"21", X"14", X"a0", X"00", X"08", 
  X"8c", X"52", X"08", X"ac", X"0f", X"f0", X"0f", X"27", 
  X"00", X"00", X"00", X"00", X"af", X"b1", X"00", X"10", 
  X"02", X"00", X"20", X"21", X"27", X"a5", X"00", X"18", 
  X"0b", X"f0", X"15", X"a7", X"00", X"00", X"30", X"21", 
  X"af", X"a5", X"00", X"28", X"0f", X"f0", X"0f", X"27", 
  X"af", X"a6", X"00", X"2c", X"8f", X"a5", X"00", X"28", 
  X"8f", X"a6", X"00", X"2c", X"af", X"b1", X"00", X"10", 
  X"02", X"00", X"20", X"21", X"02", X"40", X"f8", X"09", 
  X"00", X"40", X"38", X"21", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"3c", 
  X"24", X"03", X"00", X"8a", X"ae", X"20", X"00", X"00", 
  X"ae", X"03", X"00", X"00", X"8f", X"bf", X"00", X"3c", 
  X"8f", X"b2", X"00", X"38", X"8f", X"b1", X"00", X"34", 
  X"8f", X"b0", X"00", X"30", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"40", X"00", X"80", X"18", X"21", 
  X"3c", X"04", X"00", X"00", X"8c", X"84", X"08", X"9c", 
  X"00", X"a0", X"10", X"21", X"00", X"c0", X"38", X"21", 
  X"00", X"60", X"28", X"21", X"0b", X"f0", X"15", X"8f", 
  X"00", X"40", X"30", X"21", X"10", X"a0", X"00", X"0a", 
  X"00", X"00", X"00", X"00", X"2c", X"c2", X"01", X"00", 
  X"54", X"40", X"00", X"05", X"a0", X"a6", X"00", X"00", 
  X"24", X"02", X"00", X"8a", X"ac", X"82", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"ff", X"ff", 
  X"03", X"e0", X"00", X"08", X"24", X"02", X"00", X"01", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"27", X"bd", X"ff", X"c8", X"3c", X"02", X"00", X"00", 
  X"af", X"bf", X"00", X"34", X"af", X"b1", X"00", X"30", 
  X"af", X"b0", X"00", X"2c", X"00", X"e0", X"88", X"21", 
  X"8c", X"50", X"08", X"ac", X"af", X"a4", X"00", X"18", 
  X"af", X"a5", X"00", X"1c", X"0f", X"f0", X"0f", X"27", 
  X"af", X"a6", X"00", X"20", X"8f", X"a4", X"00", X"18", 
  X"8f", X"a5", X"00", X"1c", X"8f", X"a6", X"00", X"20", 
  X"af", X"b1", X"00", X"10", X"02", X"00", X"f8", X"09", 
  X"00", X"40", X"38", X"21", X"8f", X"bf", X"00", X"34", 
  X"8f", X"b1", X"00", X"30", X"8f", X"b0", X"00", X"2c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"38", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"00", X"80", X"88", X"21", 
  X"3c", X"10", X"00", X"00", X"00", X"a0", X"20", X"21", 
  X"00", X"c0", X"28", X"21", X"00", X"e0", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"0f", X"f0", X"06", X"58", 
  X"ae", X"00", X"0d", X"44", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"8e", X"03", X"0d", X"44", X"54", X"60", X"00", X"01", 
  X"ae", X"23", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"00", X"80", X"88", X"21", 
  X"3c", X"10", X"00", X"00", X"00", X"a0", X"20", X"21", 
  X"af", X"bf", X"00", X"1c", X"0f", X"f0", X"06", X"37", 
  X"ae", X"00", X"0d", X"44", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"8e", X"03", X"0d", X"44", X"54", X"60", X"00", X"01", 
  X"ae", X"23", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b0", X"00", X"10", 
  X"af", X"bf", X"00", X"1c", X"af", X"b2", X"00", X"18", 
  X"af", X"b1", X"00", X"14", X"14", X"a0", X"00", X"03", 
  X"00", X"a0", X"80", X"21", X"0b", X"f0", X"16", X"41", 
  X"00", X"00", X"10", X"21", X"10", X"80", X"00", X"06", 
  X"00", X"80", X"88", X"21", X"8c", X"82", X"00", X"38", 
  X"54", X"40", X"00", X"04", X"86", X"02", X"00", X"0c", 
  X"0f", X"f0", X"0b", X"91", X"00", X"00", X"00", X"00", 
  X"86", X"02", X"00", X"0c", X"10", X"40", X"00", X"25", 
  X"00", X"00", X"10", X"21", X"02", X"20", X"20", X"21", 
  X"0f", X"f0", X"0b", X"46", X"02", X"00", X"28", X"21", 
  X"00", X"40", X"90", X"21", X"8e", X"02", X"00", X"2c", 
  X"50", X"40", X"00", X"08", X"96", X"02", X"00", X"0c", 
  X"8e", X"05", X"00", X"1c", X"00", X"40", X"f8", X"09", 
  X"02", X"20", X"20", X"21", X"28", X"42", X"00", X"00", 
  X"24", X"03", X"ff", X"ff", X"00", X"62", X"90", X"0b", 
  X"96", X"02", X"00", X"0c", X"30", X"42", X"00", X"80", 
  X"50", X"40", X"00", X"05", X"8e", X"05", X"00", X"30", 
  X"8e", X"05", X"00", X"10", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"20", X"20", X"21", X"8e", X"05", X"00", X"30", 
  X"10", X"a0", X"00", X"06", X"26", X"02", X"00", X"40", 
  X"50", X"a2", X"00", X"04", X"ae", X"00", X"00", X"30", 
  X"0f", X"f0", X"0c", X"ed", X"02", X"20", X"20", X"21", 
  X"ae", X"00", X"00", X"30", X"8e", X"05", X"00", X"44", 
  X"50", X"a0", X"00", X"05", X"a6", X"00", X"00", X"0c", 
  X"0f", X"f0", X"0c", X"ed", X"02", X"20", X"20", X"21", 
  X"ae", X"00", X"00", X"44", X"a6", X"00", X"00", X"0c", 
  X"02", X"40", X"10", X"21", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b2", X"00", X"18", X"8f", X"b1", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"3c", X"02", X"00", X"00", 
  X"00", X"80", X"28", X"21", X"0b", X"f0", X"16", X"0a", 
  X"8c", X"44", X"08", X"9c", X"27", X"bd", X"ff", X"e0", 
  X"af", X"b1", X"00", X"18", X"af", X"b0", X"00", X"14", 
  X"00", X"80", X"88", X"21", X"3c", X"10", X"00", X"00", 
  X"00", X"a0", X"20", X"21", X"00", X"c0", X"28", X"21", 
  X"af", X"bf", X"00", X"1c", X"0f", X"f0", X"06", X"39", 
  X"ae", X"00", X"0d", X"44", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"8e", X"03", X"0d", X"44", X"54", X"60", X"00", X"01", 
  X"ae", X"23", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"00", X"80", X"88", X"21", 
  X"3c", X"10", X"00", X"00", X"00", X"a0", X"20", X"21", 
  X"af", X"bf", X"00", X"1c", X"0f", X"f0", X"06", X"3d", 
  X"ae", X"00", X"0d", X"44", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"8e", X"03", X"0d", X"44", X"54", X"60", X"00", X"01", 
  X"ae", X"23", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"00", X"80", X"88", X"21", 
  X"3c", X"10", X"00", X"00", X"00", X"a0", X"20", X"21", 
  X"00", X"c0", X"28", X"21", X"00", X"e0", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"0f", X"f0", X"06", X"3f", 
  X"ae", X"00", X"0d", X"44", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"8e", X"03", X"0d", X"44", X"54", X"60", X"00", X"01", 
  X"ae", X"23", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"00", X"80", X"88", X"21", 
  X"3c", X"10", X"00", X"00", X"00", X"a0", X"20", X"21", 
  X"00", X"c0", X"28", X"21", X"00", X"e0", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"0f", X"f0", X"06", X"43", 
  X"ae", X"00", X"0d", X"44", X"24", X"03", X"ff", X"ff", 
  X"14", X"43", X"00", X"05", X"8f", X"bf", X"00", X"1c", 
  X"8e", X"03", X"0d", X"44", X"54", X"60", X"00", X"01", 
  X"ae", X"23", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b0", X"00", X"14", 
  X"00", X"a0", X"80", X"21", X"8c", X"a5", X"00", X"00", 
  X"af", X"b1", X"00", X"18", X"af", X"bf", X"00", X"1c", 
  X"10", X"a0", X"00", X"03", X"00", X"80", X"88", X"21", 
  X"0f", X"f0", X"16", X"a0", X"00", X"00", X"00", X"00", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"00", X"28", X"21", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"3c", X"02", X"00", X"00", X"8c", X"42", X"08", X"9c", 
  X"27", X"bd", X"ff", X"d8", X"af", X"b0", X"00", X"14", 
  X"af", X"bf", X"00", X"24", X"af", X"b3", X"00", X"20", 
  X"af", X"b2", X"00", X"1c", X"af", X"b1", X"00", X"18", 
  X"10", X"82", X"00", X"3b", X"00", X"80", X"80", X"21", 
  X"8c", X"82", X"00", X"4c", X"00", X"00", X"88", X"21", 
  X"10", X"40", X"00", X"10", X"24", X"12", X"00", X"80", 
  X"8e", X"02", X"00", X"4c", X"00", X"51", X"10", X"21", 
  X"8c", X"45", X"00", X"00", X"50", X"a0", X"00", X"06", 
  X"26", X"31", X"00", X"04", X"8c", X"b3", X"00", X"00", 
  X"0f", X"f0", X"0c", X"ed", X"02", X"00", X"20", X"21", 
  X"0b", X"f0", X"16", X"c3", X"02", X"60", X"28", X"21", 
  X"56", X"32", X"ff", X"f6", X"8e", X"02", X"00", X"4c", 
  X"8e", X"05", X"00", X"4c", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"00", X"20", X"21", X"8e", X"05", X"00", X"40", 
  X"50", X"a0", X"00", X"04", X"8e", X"05", X"01", X"48", 
  X"0f", X"f0", X"0c", X"ed", X"02", X"00", X"20", X"21", 
  X"8e", X"05", X"01", X"48", X"54", X"a0", X"00", X"08", 
  X"26", X"12", X"01", X"4c", X"8e", X"05", X"00", X"54", 
  X"50", X"a0", X"00", X"0e", X"8e", X"02", X"00", X"38", 
  X"0f", X"f0", X"0c", X"ed", X"02", X"00", X"20", X"21", 
  X"0b", X"f0", X"16", X"e7", X"8e", X"02", X"00", X"38", 
  X"50", X"b2", X"ff", X"f9", X"8e", X"05", X"00", X"54", 
  X"8c", X"b1", X"00", X"00", X"0f", X"f0", X"0c", X"ed", 
  X"02", X"00", X"20", X"21", X"12", X"32", X"ff", X"f3", 
  X"02", X"20", X"28", X"21", X"0b", X"f0", X"16", X"e1", 
  X"8c", X"b1", X"00", X"00", X"10", X"40", X"00", X"0f", 
  X"8f", X"bf", X"00", X"24", X"8e", X"02", X"00", X"3c", 
  X"00", X"40", X"f8", X"09", X"02", X"00", X"20", X"21", 
  X"8e", X"05", X"02", X"e0", X"10", X"a0", X"00", X"08", 
  X"8f", X"bf", X"00", X"24", X"8f", X"b3", X"00", X"20", 
  X"8f", X"b2", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"02", X"00", X"20", X"21", X"8f", X"b0", X"00", X"14", 
  X"0b", X"f0", X"16", X"a0", X"27", X"bd", X"00", X"28", 
  X"8f", X"bf", X"00", X"24", X"8f", X"b3", X"00", X"20", 
  X"8f", X"b2", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"3c", X"04", X"bf", X"c0", 
  X"27", X"bd", X"ff", X"e8", X"af", X"bf", X"00", X"14", 
  X"0f", X"f0", X"06", X"66", X"24", X"84", X"5c", X"60", 
  X"3c", X"04", X"bf", X"c0", X"0f", X"f0", X"06", X"66", 
  X"24", X"84", X"5c", X"70", X"3c", X"04", X"bf", X"c0", 
  X"0f", X"f0", X"06", X"8a", X"24", X"84", X"5c", X"98", 
  X"3c", X"04", X"bf", X"c0", X"24", X"84", X"5c", X"b0", 
  X"0f", X"f0", X"06", X"8a", X"24", X"05", X"00", X"2a", 
  X"8f", X"bf", X"00", X"14", X"00", X"00", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"18", 
  X"30", X"30", X"30", X"30", X"30", X"30", X"30", X"30", 
  X"30", X"30", X"30", X"30", X"30", X"30", X"30", X"30", 
  X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
  X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
  X"0a", X"0a", X"4c", X"69", X"62", X"43", X"20", X"54", 
  X"65", X"73", X"74", X"0a", X"00", X"00", X"00", X"00", 
  X"63", X"6f", X"6d", X"70", X"69", X"6c", X"65", X"20", 
  X"74", X"69", X"6d", X"65", X"3a", X"20", X"46", X"65", 
  X"62", X"20", X"32", X"30", X"20", X"32", X"30", X"31", 
  X"34", X"20", X"2d", X"2d", X"20", X"32", X"30", X"3a", 
  X"35", X"30", X"3a", X"33", X"32", X"00", X"00", X"00", 
  X"67", X"63", X"63", X"20", X"76", X"65", X"72", X"73", 
  X"69", X"6f", X"6e", X"3a", X"20", X"20", X"34", X"2e", 
  X"38", X"2e", X"31", X"0a", X"00", X"00", X"00", X"00", 
  X"0a", X"0a", X"54", X"68", X"69", X"73", X"20", X"69", 
  X"73", X"20", X"61", X"20", X"70", X"72", X"69", X"6e", 
  X"74", X"66", X"20", X"74", X"65", X"73", X"74", X"3a", 
  X"20", X"25", X"64", X"0a", X"0a", X"00", X"00", X"00", 
  X"30", X"31", X"32", X"33", X"34", X"35", X"36", X"37", 
  X"38", X"39", X"41", X"42", X"43", X"44", X"45", X"46", 
  X"00", X"00", X"00", X"00", X"30", X"31", X"32", X"33", 
  X"34", X"35", X"36", X"37", X"38", X"39", X"61", X"62", 
  X"63", X"64", X"65", X"66", X"00", X"00", X"00", X"00", 
  X"43", X"00", X"00", X"00", X"50", X"4f", X"53", X"49", 
  X"58", X"00", X"00", X"00", X"2e", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"02", X"ec", 
  X"00", X"00", X"03", X"50", X"00", X"00", X"03", X"b4", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"bf", X"c0", X"5c", X"f8", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", 
  X"33", X"0e", X"ab", X"cd", X"12", X"34", X"e6", X"6d", 
  X"de", X"ec", X"00", X"05", X"00", X"0b", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"41", X"53", X"43", X"49", X"49", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"41", X"53", X"43", X"49", X"49", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"bf", X"c0", X"5d", X"04", X"bf", X"c0", X"5c", X"ac", 
  X"bf", X"c0", X"5c", X"ac", X"bf", X"c0", X"5c", X"ac", 
  X"bf", X"c0", X"5c", X"ac", X"bf", X"c0", X"5c", X"ac", 
  X"bf", X"c0", X"5c", X"ac", X"bf", X"c0", X"5c", X"ac", 
  X"bf", X"c0", X"5c", X"ac", X"bf", X"c0", X"5c", X"ac", 
  X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", 
  X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"04", X"90", X"00", X"00", X"04", X"90", 
  X"00", X"00", X"04", X"98", X"00", X"00", X"04", X"98", 
  X"00", X"00", X"04", X"a0", X"00", X"00", X"04", X"a0", 
  X"00", X"00", X"04", X"a8", X"00", X"00", X"04", X"a8", 
  X"00", X"00", X"04", X"b0", X"00", X"00", X"04", X"b0", 
  X"00", X"00", X"04", X"b8", X"00", X"00", X"04", X"b8", 
  X"00", X"00", X"04", X"c0", X"00", X"00", X"04", X"c0", 
  X"00", X"00", X"04", X"c8", X"00", X"00", X"04", X"c8", 
  X"00", X"00", X"04", X"d0", X"00", X"00", X"04", X"d0", 
  X"00", X"00", X"04", X"d8", X"00", X"00", X"04", X"d8", 
  X"00", X"00", X"04", X"e0", X"00", X"00", X"04", X"e0", 
  X"00", X"00", X"04", X"e8", X"00", X"00", X"04", X"e8", 
  X"00", X"00", X"04", X"f0", X"00", X"00", X"04", X"f0", 
  X"00", X"00", X"04", X"f8", X"00", X"00", X"04", X"f8", 
  X"00", X"00", X"05", X"00", X"00", X"00", X"05", X"00", 
  X"00", X"00", X"05", X"08", X"00", X"00", X"05", X"08", 
  X"00", X"00", X"05", X"10", X"00", X"00", X"05", X"10", 
  X"00", X"00", X"05", X"18", X"00", X"00", X"05", X"18", 
  X"00", X"00", X"05", X"20", X"00", X"00", X"05", X"20", 
  X"00", X"00", X"05", X"28", X"00", X"00", X"05", X"28", 
  X"00", X"00", X"05", X"30", X"00", X"00", X"05", X"30", 
  X"00", X"00", X"05", X"38", X"00", X"00", X"05", X"38", 
  X"00", X"00", X"05", X"40", X"00", X"00", X"05", X"40", 
  X"00", X"00", X"05", X"48", X"00", X"00", X"05", X"48", 
  X"00", X"00", X"05", X"50", X"00", X"00", X"05", X"50", 
  X"00", X"00", X"05", X"58", X"00", X"00", X"05", X"58", 
  X"00", X"00", X"05", X"60", X"00", X"00", X"05", X"60", 
  X"00", X"00", X"05", X"68", X"00", X"00", X"05", X"68", 
  X"00", X"00", X"05", X"70", X"00", X"00", X"05", X"70", 
  X"00", X"00", X"05", X"78", X"00", X"00", X"05", X"78", 
  X"00", X"00", X"05", X"80", X"00", X"00", X"05", X"80", 
  X"00", X"00", X"05", X"88", X"00", X"00", X"05", X"88", 
  X"00", X"00", X"05", X"90", X"00", X"00", X"05", X"90", 
  X"00", X"00", X"05", X"98", X"00", X"00", X"05", X"98", 
  X"00", X"00", X"05", X"a0", X"00", X"00", X"05", X"a0", 
  X"00", X"00", X"05", X"a8", X"00", X"00", X"05", X"a8", 
  X"00", X"00", X"05", X"b0", X"00", X"00", X"05", X"b0", 
  X"00", X"00", X"05", X"b8", X"00", X"00", X"05", X"b8", 
  X"00", X"00", X"05", X"c0", X"00", X"00", X"05", X"c0", 
  X"00", X"00", X"05", X"c8", X"00", X"00", X"05", X"c8", 
  X"00", X"00", X"05", X"d0", X"00", X"00", X"05", X"d0", 
  X"00", X"00", X"05", X"d8", X"00", X"00", X"05", X"d8", 
  X"00", X"00", X"05", X"e0", X"00", X"00", X"05", X"e0", 
  X"00", X"00", X"05", X"e8", X"00", X"00", X"05", X"e8", 
  X"00", X"00", X"05", X"f0", X"00", X"00", X"05", X"f0", 
  X"00", X"00", X"05", X"f8", X"00", X"00", X"05", X"f8", 
  X"00", X"00", X"06", X"00", X"00", X"00", X"06", X"00", 
  X"00", X"00", X"06", X"08", X"00", X"00", X"06", X"08", 
  X"00", X"00", X"06", X"10", X"00", X"00", X"06", X"10", 
  X"00", X"00", X"06", X"18", X"00", X"00", X"06", X"18", 
  X"00", X"00", X"06", X"20", X"00", X"00", X"06", X"20", 
  X"00", X"00", X"06", X"28", X"00", X"00", X"06", X"28", 
  X"00", X"00", X"06", X"30", X"00", X"00", X"06", X"30", 
  X"00", X"00", X"06", X"38", X"00", X"00", X"06", X"38", 
  X"00", X"00", X"06", X"40", X"00", X"00", X"06", X"40", 
  X"00", X"00", X"06", X"48", X"00", X"00", X"06", X"48", 
  X"00", X"00", X"06", X"50", X"00", X"00", X"06", X"50", 
  X"00", X"00", X"06", X"58", X"00", X"00", X"06", X"58", 
  X"00", X"00", X"06", X"60", X"00", X"00", X"06", X"60", 
  X"00", X"00", X"06", X"68", X"00", X"00", X"06", X"68", 
  X"00", X"00", X"06", X"70", X"00", X"00", X"06", X"70", 
  X"00", X"00", X"06", X"78", X"00", X"00", X"06", X"78", 
  X"00", X"00", X"06", X"80", X"00", X"00", X"06", X"80", 
  X"00", X"00", X"06", X"88", X"00", X"00", X"06", X"88", 
  X"00", X"00", X"06", X"90", X"00", X"00", X"06", X"90", 
  X"00", X"00", X"06", X"98", X"00", X"00", X"06", X"98", 
  X"00", X"00", X"06", X"a0", X"00", X"00", X"06", X"a0", 
  X"00", X"00", X"06", X"a8", X"00", X"00", X"06", X"a8", 
  X"00", X"00", X"06", X"b0", X"00", X"00", X"06", X"b0", 
  X"00", X"00", X"06", X"b8", X"00", X"00", X"06", X"b8", 
  X"00", X"00", X"06", X"c0", X"00", X"00", X"06", X"c0", 
  X"00", X"00", X"06", X"c8", X"00", X"00", X"06", X"c8", 
  X"00", X"00", X"06", X"d0", X"00", X"00", X"06", X"d0", 
  X"00", X"00", X"06", X"d8", X"00", X"00", X"06", X"d8", 
  X"00", X"00", X"06", X"e0", X"00", X"00", X"06", X"e0", 
  X"00", X"00", X"06", X"e8", X"00", X"00", X"06", X"e8", 
  X"00", X"00", X"06", X"f0", X"00", X"00", X"06", X"f0", 
  X"00", X"00", X"06", X"f8", X"00", X"00", X"06", X"f8", 
  X"00", X"00", X"07", X"00", X"00", X"00", X"07", X"00", 
  X"00", X"00", X"07", X"08", X"00", X"00", X"07", X"08", 
  X"00", X"00", X"07", X"10", X"00", X"00", X"07", X"10", 
  X"00", X"00", X"07", X"18", X"00", X"00", X"07", X"18", 
  X"00", X"00", X"07", X"20", X"00", X"00", X"07", X"20", 
  X"00", X"00", X"07", X"28", X"00", X"00", X"07", X"28", 
  X"00", X"00", X"07", X"30", X"00", X"00", X"07", X"30", 
  X"00", X"00", X"07", X"38", X"00", X"00", X"07", X"38", 
  X"00", X"00", X"07", X"40", X"00", X"00", X"07", X"40", 
  X"00", X"00", X"07", X"48", X"00", X"00", X"07", X"48", 
  X"00", X"00", X"07", X"50", X"00", X"00", X"07", X"50", 
  X"00", X"00", X"07", X"58", X"00", X"00", X"07", X"58", 
  X"00", X"00", X"07", X"60", X"00", X"00", X"07", X"60", 
  X"00", X"00", X"07", X"68", X"00", X"00", X"07", X"68", 
  X"00", X"00", X"07", X"70", X"00", X"00", X"07", X"70", 
  X"00", X"00", X"07", X"78", X"00", X"00", X"07", X"78", 
  X"00", X"00", X"07", X"80", X"00", X"00", X"07", X"80", 
  X"00", X"00", X"07", X"88", X"00", X"00", X"07", X"88", 
  X"00", X"00", X"07", X"90", X"00", X"00", X"07", X"90", 
  X"00", X"00", X"07", X"98", X"00", X"00", X"07", X"98", 
  X"00", X"00", X"07", X"a0", X"00", X"00", X"07", X"a0", 
  X"00", X"00", X"07", X"a8", X"00", X"00", X"07", X"a8", 
  X"00", X"00", X"07", X"b0", X"00", X"00", X"07", X"b0", 
  X"00", X"00", X"07", X"b8", X"00", X"00", X"07", X"b8", 
  X"00", X"00", X"07", X"c0", X"00", X"00", X"07", X"c0", 
  X"00", X"00", X"07", X"c8", X"00", X"00", X"07", X"c8", 
  X"00", X"00", X"07", X"d0", X"00", X"00", X"07", X"d0", 
  X"00", X"00", X"07", X"d8", X"00", X"00", X"07", X"d8", 
  X"00", X"00", X"07", X"e0", X"00", X"00", X"07", X"e0", 
  X"00", X"00", X"07", X"e8", X"00", X"00", X"07", X"e8", 
  X"00", X"00", X"07", X"f0", X"00", X"00", X"07", X"f0", 
  X"00", X"00", X"07", X"f8", X"00", X"00", X"07", X"f8", 
  X"00", X"00", X"08", X"00", X"00", X"00", X"08", X"00", 
  X"00", X"00", X"08", X"08", X"00", X"00", X"08", X"08", 
  X"00", X"00", X"08", X"10", X"00", X"00", X"08", X"10", 
  X"00", X"00", X"08", X"18", X"00", X"00", X"08", X"18", 
  X"00", X"00", X"08", X"20", X"00", X"00", X"08", X"20", 
  X"00", X"00", X"08", X"28", X"00", X"00", X"08", X"28", 
  X"00", X"00", X"08", X"30", X"00", X"00", X"08", X"30", 
  X"00", X"00", X"08", X"38", X"00", X"00", X"08", X"38", 
  X"00", X"00", X"08", X"40", X"00", X"00", X"08", X"40", 
  X"00", X"00", X"08", X"48", X"00", X"00", X"08", X"48", 
  X"00", X"00", X"08", X"50", X"00", X"00", X"08", X"50", 
  X"00", X"00", X"08", X"58", X"00", X"00", X"08", X"58", 
  X"00", X"00", X"08", X"60", X"00", X"00", X"08", X"60", 
  X"00", X"00", X"08", X"68", X"00", X"00", X"08", X"68", 
  X"00", X"00", X"08", X"70", X"00", X"00", X"08", X"70", 
  X"00", X"00", X"08", X"78", X"00", X"00", X"08", X"78", 
  X"00", X"00", X"08", X"80", X"00", X"00", X"08", X"80", 
  X"00", X"00", X"08", X"88", X"00", X"00", X"08", X"88", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"01", X"ff", X"ff", X"ff", X"ff", 
  X"00", X"02", X"00", X"00", X"bf", X"c0", X"56", X"f4" 
  );

constant INIT_DATA : t_obj_code(0 to 199) := (
  X"30", X"30", X"30", X"30", X"30", X"30", X"30", X"30", 
  X"30", X"30", X"30", X"30", X"30", X"30", X"30", X"30", 
  X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
  X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
  X"0a", X"0a", X"4c", X"69", X"62", X"43", X"20", X"54", 
  X"65", X"73", X"74", X"0a", X"00", X"00", X"00", X"00", 
  X"63", X"6f", X"6d", X"70", X"69", X"6c", X"65", X"20", 
  X"74", X"69", X"6d", X"65", X"3a", X"20", X"46", X"65", 
  X"62", X"20", X"32", X"30", X"20", X"32", X"30", X"31", 
  X"34", X"20", X"2d", X"2d", X"20", X"32", X"30", X"3a", 
  X"35", X"30", X"3a", X"33", X"32", X"00", X"00", X"00", 
  X"67", X"63", X"63", X"20", X"76", X"65", X"72", X"73", 
  X"69", X"6f", X"6e", X"3a", X"20", X"20", X"34", X"2e", 
  X"38", X"2e", X"31", X"0a", X"00", X"00", X"00", X"00", 
  X"0a", X"0a", X"54", X"68", X"69", X"73", X"20", X"69", 
  X"73", X"20", X"61", X"20", X"70", X"72", X"69", X"6e", 
  X"74", X"66", X"20", X"74", X"65", X"73", X"74", X"3a", 
  X"20", X"25", X"64", X"0a", X"0a", X"00", X"00", X"00", 
  X"30", X"31", X"32", X"33", X"34", X"35", X"36", X"37", 
  X"38", X"39", X"41", X"42", X"43", X"44", X"45", X"46", 
  X"00", X"00", X"00", X"00", X"30", X"31", X"32", X"33", 
  X"34", X"35", X"36", X"37", X"38", X"39", X"61", X"62", 
  X"63", X"64", X"65", X"66", X"00", X"00", X"00", X"00", 
  X"43", X"00", X"00", X"00", X"50", X"4f", X"53", X"49", 
  X"58", X"00", X"00", X"00", X"2e", X"00", X"00", X"00" 
  );



end package OBJ_CODE_PKG;
